`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
DeGy5rZwNuOJnxDZjckajf3bMqwWif4RCyd05MX0eywgMTnKoLl1RONDF4yQFeTIkRdBucpGR1iq
WAwTqzDsgw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Ielrw6BZF3pVyiPC9RrKbpA6zsA//x1ypIetoDu5OLW185egTvFvEaSvEavdXIyvJ6TqtQ50Zy07
i+XVo2hi9kgmV1dUe0hFouhINyHywDQ0CAGTpeqGRqWGZ51ri8DbgyTG5wnHVxFah6s+/bLrxhFl
M/+AMw+v4ENWezwbMVo=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Lk+Q58K/N2QIcYtYIKwe6ta5UtwJ70247eA1ClsuIXDa2pu7qmuCX51/DpdSJTW/Jusfwa69lYFb
GBfXNtjiUOMa0Qe5e+ofgi1ySq/SyQUIFM8R8ftVQ+OxqjSO/CslAjUkekGqBS2ltjDEGnMqvLAo
M7sSOHTYK/tgudKAthR3MYZNVocUufH47B6tiZxrjADqo+yI71wi7Cmdq5u0NFa5Rxm5QMxQm5u2
mYhbObMpii8qPjGUKmvFU4TJmeH8f+JZcGCIYwSNIgh/kgMiDPz7xR/fNtpm4WfoREjxYV+d2MjR
3DMNd5N8VVYkGYzK6DQHD7xHShwg8t1+Y+ZzSg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
W0oMsx7XqXE7ZbjkkRdJD1BDlVkUJsSw3N7P8Y2rwpp7a+/6kgYjXXrNLBKeb81kYMtWqxwtqGlU
WDIqIEoIW1muxnFT92jKGo69ZkBhq4qB4VmPU/ppb4mC8MGtDikzxGCrIYHNnJN0LoH5bldVtL5P
6PAcA58bm92Qb2MoC3McU/oACY86Pd8gS72PUtj5SwxyQQ9X4z6Z9x8wf8kfNMLQQkhpnmmwcTBY
JBTnne+vE7hGOyedXEA+8Iymy7yKHiWJF3Eihf64wNlQd8O14ejMwDbbm+QRwmcz541Le/7wkXJy
t0s8Vk+Lyd48uolBljYcYuesqEm7ZamuacXcdg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
tQ81J0IMscjxt9p9FIkV7dqh9WgOclKcyzlSCz98RRq+PVggE0ECzkxdaoh/0Sl44A9lH0VOOsCr
crHiz2R3lXz7OI7uoYSuOeVhLAkJgJ3w6//ArWvrIPnIc/BEKopj27R4cfmtD9KDBKnFctiY4CWZ
M3SDuVFIBlElwo8PCdosvm19J5sO1NeuRmgsQOtylQiiGFyE7wgPV1HvXOJ8tkMlr1oKS7SRlyVQ
R9ux1BJhOOvkzoFctKzAAtb1rKgXwb9Kv/aGh2rgGL5bQBh7oNqCNo/YeYYExeetQfZLXtda9nmr
Iu3gvXKYLDl4PJt+PyzqmrE5htCyBjcA1FZjjw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
mTvyfHTcYgSTrB9qQYYZTd5LTrftm8mzmwAYim4QlJecmM0jwEIRJdrI02IKhoHDRp4is1o0feqc
bZgTDyGWdny3SkOXfQG7L+LRfWZhhEsFrOAeD/ognlNQeEvO1qy17GxJ6MNHZ3vY6T1xMtEv6SC6
mWMFT6G55O8/Ocylhgc=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
T7ekYXsF8w6cT4y8Sp1k0Ytg9aQzWDsMR4Q2RkSkokYPmbvJfUOCpmYDknFj5pXzlRBxFioxZVGk
julh1nbAoh7oAXXxhF/WDpVTggOqJNBAOBXqix2rLR/x/CKnxo0fLnsJChIaisJUsr0aRsMUlMW8
ehbQeFodvLjulg4EEW2qD9fYeMC3DTi9n8sV2zk1UNmAcmsW7JQeqDtkPZmNiovvDd7Vv23I8ePj
tBprvHFzz/27ATNB5Z4+toWCXik5Du0udlT8plpo+FlKlqafgSgJqERthq6folUni3c09aq8e2H0
FS8CZq7zJg/ncBQCJVZWqfjzKSgDLQ47F/b2yw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15104)
`pragma protect data_block
MScHo31tlAUz550tzvz8yqM6U63qUR1DQGqR+LSK284rtYjdqVgER10Agik+kE5hHBCXX7Sqi96P
e7V2CfT0jtbpMMpTlfAJg8ZfuNfGaj2SEONykZyLc8yo19R5sgSJUd/Si81fgGXxZAJp1di5FQ98
n/Vt+spqloYdulUwZgXvDF6zQQFrpiCITWIlJ8ktwxGLPPD0XkGtQMsR/q8fW5SDw31FUnl9LVE3
KWDxAbDyZW8VRRI3cnon0MYLNIoH1FNjQ/0hkJNTlp4RfP9cp8Ae5cgKekwEeeQRmDW5xtUMH6xN
4T6TfsxAlLpXGdEWVj6/gBSu5ZtHbHrv9tRGehI7bSPoVupAQ6+bmvjIbqWFKsFm7xrYOn9Vl9g+
R7vy4aACynPJ3b7wxIaqZlFzLp31MVB/RthtgRFLUq2aGU5l5Hfdnb4upkzgVUsmQpYcEVaiz16s
DIcQeXJOL/EnjgFniwTiaHp+wnc8sZt4O3EalON/0lnUak6hTsaJ2xd31X8YWraTpxdw9QglFAdW
JhJnEVetHFyK25qpundbAMMaZKGyXPAFi57mnrzQ4tJvympCwFinXhTkuYxiu8VON+dDyVs7VxWt
mll7Nr8IO4CoGcelXe0RpI+x8B+c80W1bLgTtISgbMBo1xf8b1iQdAkcZwVbGS9AOHzEDNIycLdm
tXnNu/e/I6Zn+0bMYAUPw80XSS7rZc6b4xCZ3aiugiRPNVvWprmJ2ePBDURNx34yDckSEWfXYZsJ
RffaJMK0S2/NfYabvWPT14uZpekG0AiNfTwfXTvFOwbXPmoLbDNy1/UAZOGl4VNX9+sDaL5f7qTd
SN7ryjDvZfX9+mH9GRBI2mHJaYw7GUXcSssqWwXPp8XYqgMER0ijllzyhlw1L9KaxpHM1oH4pcT9
7hhh96YzgcOnzYxfD4ORyXpxj8JSMWoaEdoLZF7OLR2AXbJU1jXV+xl11x9jNYHl8BURWQtRAEYD
0dUmcX4M0lQ1wcEezBQOyfXzZaFFeWL9ZRWX0l26AK4Pj1sd4rZw26dXbI6NMQ7sgdJ1NTLMUVYk
u+Mw7knW/StoBkqChJztvgHC7OcsdDq1oUcB10+syHHCh6G2QQQQ9F3Gx4H/LVTOqy/au/FOk0SC
tQN10QCDCQJhBHAfpxyOjWz1vWf2kglIgGzC3iAuKH+41cmxLWg93wqVKjax5cbVDklATs1L0zJ5
kqjP6C6DllcYUeIDh9l5v9/i4+U/5Y0ZdAwEsLfIQLFKaRNOm5oSNMOOeGEYBiXegzcFZsq/lw7n
aDhh7pCV2TkLsXhYx5wLoGBToAaWQtzmGOuWoBS3ay+CqwzVhztHs0lWTF1M10VgT183CbrfXVGb
CSZBKiCvOrRB/ZrZPH+VRDu910gzQGbBnRQjUwc527U4rDMjVsgAxKWTnc6BXnvyLr3ZxtZiQvMY
LrXwL6RBWLXZiqWjDoyHGWlPai7nRvkyoH8zP4JRGYy+nzCmvaDnvzCnjN4AI6sTr0fUIiOd9Sz/
4becsjsUuwSmyvbmuPOOZ3itPoVO10c6Uhy/swI4dDJdQ9B4dlmu7BeOSb0m7tFyHpUzqxWlKXUx
wPBUWZRgpDspeYZ4jc6hHzfiYNqFd1VMYkD2r8ArkSyKCmj6N+36BcDFXYyNtySK/LtF31mQfkW5
SL2Xue9fsuglEZSYJrTEMak21fn30Ektzw9i5ynFSEdxKRNgticD95lFt9CVQdQw9E91qwpVGmhz
bBafGT3CbaGGTmfuxH+wta5bfn4bBuW+ZAVp6VAIIoRljKHfPQ6xTN4KI0dq8qz5SqtQiRhk6DVh
b0i6wk0ehtucVxKUX0221Zqj70MprLhFxNhNyWb5n7ueQFIU6IbRfS6n2ehuv7wAJqxoDeY9IqM1
ysK+d6/oE15YSSghzSMWN+cUIzlJ80DxvDUVcYm9VbkvA1eBXqquM4ud116WvfpAZokciI4GzaW2
gytNuhdgY9iWoGRODdg2n4i6j0QqmK/8eLbkLB1oRDbGIZgUTyXadoRTKgX1eAtrgcgkj9LfkSI3
7/vcSY02nAb0nPZsOUbXx9lNu/lvCoCsDEJVrxoDgwd7kYCGzNK62ukvA36N9ptjgo7Sh1AMlyxo
Na0/r7tXliwalifKCkoU8SnK1SLPMBkEdDaXbju4lRW4ibVCqZe4SUcYRWlJ84Tty/OKqK/PmTfq
15ByUiyY+2POYTCtNBPG1050NA802rAtc998FDcp4yoY9jBvvVD5pljMiPeliBV2MMTz8pXX14Nr
koeKMiUobIxioaof/loLzZ7vkfpgsLyKpWv76u/6krdAQ2ABBLjgRGaYhfVMeaiJJES5K1/HXONz
2bKeJCCk7p16wZ5/x1W+yFqjnohczLX39buscFWPD2sWxp9nQTUxg59CbaToB0WwL3g8zwp0ULHM
lDYuqiz+8LKgZvCm5fT2TMTmsMnD1eJWob9apiK3lrYCKsr0I6WDkU6bfshiK2NSF9yXhrN7nTr/
6JRY7i74+9Pcz44s+ren3itEfhi2vqj8+dUugCHr7tvfH2671w9JqWvoLJkN1/5GsOXoLfW9/wOT
j/Y+nw6j1PGc7yo8vs96FetYGd1YCdFRDbF3WNddMCRdvm+ZvjVPYAIJBSzhjAXJB7zXd3x5v7T/
GC/hs/YvYQ8wEACcWNplMtBFP3wWOX6dAGxAj46r6JghEJ11H/nnekLaUMPVQGrWnTOepWMRXSdj
OsKUF1UUxGSkwlCK5nhv9rfrIjLho3evD7G6P5wgYlnKy+l5kcX73tdoEsXWgSGdy24tkrxikCak
5RaxTs8Arr7uKfiQ4lJG+MBHOKbHava01VP8aKXzwar0so4w6sLJ7vdJsF2jqkBG5potf+di5SWg
VztusdoZiVLx9Xs0JwJufWqmPPdQryUuOjZrotp+KJLnbu99PpwEh4H1XxyCrvIkQNo9kXYBrAdx
sT+hJyr0BWryTMOt37XWzS8oy/TELhAU8MvfkDE32LX3DrviJtfo3MOTL724P62bBqUjNHYVR9ui
SW+WifM+A0KHsf95i61yPKTV4hXjtepNAgNdjsO1gXhpvfVhet/ZxcuAjUjbhNLKDZ9Cd1t6N2iS
sJPETZtJ3MkP5QvkifPHDm4YzTEmripK7ULGU5uLxBsPgyn5gwfnq14U/dCW98itoqLNuiEZjUrH
nRX9ryJmC7xawmSlLqSj03o6VpkhroY0ptM+MyN/KB4ktk45w/XgeJVbHrInPJvTd1GY3Elouxno
3B7smlPS0vQxPIL6idSosGSmKOwhjiF5oNKVGmGC3yBGNkD5b1UaQ7r+kZniKUvYnVFkcgTJBrwE
QvQyy9FoDQPlsit/xoYRoRhGlG4kXn3rktG116dd+EAaMZw/6mk2dz3quH1sKQhSt8JavnPyKV6u
WfwXJKuiktHsmunXbKBKKQ7hvcWsPBNgteJx2cRYMrItinyC+sihMjRImITANZOCQ5NnIiMM2G7o
G0cghnby/tpHrJxixcQU2sIkyOy9tcj8z4EwoBS4KHbQ6TDQ7zy17QEIwMtiHdj6aYCwnK41Im5Y
04Q1F8OsB1+TAKIHBHZcx1D2ARzsNCrq2/DlYNXWvDlACIZWx36LKZNwi2qszB4J97b7ORKzRoVh
/RZwEvIY9vAuGM3X5J1o2U97mOBiT77Sjew5LAcdS2v6CFsYw2P92DT+ghtELXnDdcFIUu48mmo4
H0p+E/h/R9BLOdgqvp3iABV6EyeABAfqkVAt9q58OZfCeIfFPRxo2+yuByKzAoCDCClopX7/OE49
l8fOVG/6y3BXbxhBs/HtT1p6AZOD8HVOsXvbs6iuuhLbHtjCwrt8FdRfAsKK0Dq/525xb2/SBQvm
vZyyl2L0O8xTQjwqzuwfVL/MKwo131g5TQfenwqQFsLUc8vcbhxK67Aniei42rbrOzMVh0KnIKNC
S0vOQv2aSmiEtXUCQLTG9h6/Cpkn4sj90/K+xiS+wB74Jkyija7HUQAKXSyiXX3qSo2OekylsPO3
1jP0G53QaCnMue0JVlj66ZZEUEpwDum9ZM9i1FYuFoHT64qgo0NTrDTLb89oBMKwuU5rSFohzmLb
o/CRdQ1BrDg6tCjKGWVBQxFDAOyeyqTxIAde7wXwfdywBGH/UG53AHo1zlVzkt/wMydcQoqYIipv
iRnDszNVAGN8nzW3WnqNMmu6kJbIzPWjiaeaarSkGOHElwESHAxs1G1+SNq3U+Hd3AfLIj1sv5Gf
CMEhg/n/GMBDyYG+nLC6NPQEq7MqqUJai0X4QZPbZjP/NZ/9kQO5DlMdU5doFAHarPINTqD0W2AD
Oiz+2lSB8Jgh5S5Lj+mMDnMje7vN0KDTdZwIeB3+30dHVxgOwof3JQtMJnvs7kHGIIFxuMwIhjBj
8ikxATcstEuikJ1td7UFJ/k+oPjIMCTRTq2huVhHZHOUR6ICdAUthoivxoMwPKcj0PpGtByDyB9o
nyfDL/QgTvnithuNDeuUJc7zOFG7KJAxP46M/Vrt58p7m+yg0SCBVpdX2IknlQEGabJyXtFMZ6U5
HUhh2hI7J4Bm6BIqD5+yMzCLfcfdWkqIMkl2Qfkuj6fKqVcY6YBr35sEfQLrYhxoYAaOp2UlDlba
wr3up3/AhFh8dg24CyPwozHdlq9pV8j8PNgjLl7YBT9TuyFf2uNVMtJ6+q5ctbuxfix+r0P5IMdL
XyOA3IOoQcsHJSyj1B+CJpbc8DFh7FhgbgwW1MxjBXGbad+PglcJoJ5nkQc91Pbzmstjh9Wiyb3M
OTroidD/hoGJYLg0ddZdRGiTjqzLSa6NkXn3sg6oTQpcFtSU84T73V3fEQsg8veQdCNqKpRX75/7
crnzI/T46F5qaj3+E3bMh8tfqb8m/XOYAp4wJMv8aGl05mkO3mpw4+O+ImIUytdiRClShnJpfrov
Zu3qZTrSaTknUI/dSPvLvPnZW/z4iQEdqrEQ77k7NW9yVwIblzhh/PWY6aPpOBt2qUM9Qwv1Ezi7
E+nIMmFa8v8sXWNA/s71rARPJUEMx22yzamlD8PurLW8DbnqCEh42YQZ5F3OFPuGALsj7Rzleqc+
cGipE9SVoLu31OlTMpDf7T/5WvH+bPysp4KAxZVUjMp6HhljOTtxT6oDaWV7XCCYVU94Cchrm/jG
5xVibst39y0x940tkHus3hti2x5UQ48O2nGKPlg7cz3SPqQ4bTxXsbxtr9CcBpiPi/+1QptEHf1p
kjnSsJdGKKmfYQ6Q2cdRyB3ZzMwNjZcUeBPdWKOgOkBJKdmdUqL5rE74qLlgKrA071zS+mEBFk1c
VU4JeHLM5Zobr9Jj1+ma01nIDEPYCHB3NpDv16YCTq0HB17nT+ITjt06EnwzXg6nDnMjn7A4Zj7v
vj5lWnVc4xlkxzv7HCn1WZQf2xojLMallngE5hefX/eWfnpolQPF3JzprjFVHDJ721xJ/1rU4ywH
waH25uilNDyxJASYtpnN7swWodsB1U2vCt/pUJvxIicl0xxoz5Iyg5jVErAyqJG65cnkAS//1QoF
IGq3SQ68rsZbOlTIcX6NDoR7F/OZscfzyJOh4nYK1QIXPvo+RuT9GgiSuCVI2z98yn/NjSHGMyD6
2WPEbM1crHWhTB03Bi5wETjZOT2c3zb6u7qfYiYmqAVQmHtb9V1eNce4DxlLNQYYdiNTMg6wUMTE
YO2uj1QoB3SujU/kCHBz4HLDqI2L1qpamKEebnObKpAFzMH1/P+F7pwBJvHU8MyCGH4NfH8GTDfS
Bxc+6Bk8wGaEVRmS04ibJyCXlw23sySm+JMHl26kQ0OCz88O3z1KiKpXXoZlVABA//dCpcD9FFpv
YWYiWdv9KB323TuDb6OXK7+/NqLBe+f/r01F4zNoW4o+iJlwD79B8TIhaeRi98gQfPOrVRDscifF
JjEVz9IXR5uQQBeB//gbBqqZWESTVKI8AEsIUwxvoGqXHx+HM3bQmVZxdkLfm1KvqmwShiuVgHuE
GPbgNf0fNlsSATEtsofitZRBF1UkNDSZek0KgvO8yuo16wTzcW8sXyBJDCzSXUiOf94BG6hQnmBs
+2yeAVD6XepwjPZnfE5cHVl3XwH7j6D7az/tid0reg+OTF7VXd9m3gyVxFHGk/h3cDj14CktOwgk
PtebPQ52q2eZ9r+8TT6GX4zsa68sJcu9BkEJnTLyr2Rfx4HyaLJqIEbIBp0Cqs8qftkB7ok7X6KJ
Zb7C7lCSMWgQNNKqCjuOSJwID4IhVNsGfrztAO+sGtOSKsbj/K05rcr2rwCDES0LBjK35w5wYeBT
c+mquoYFdYYkqyvCJrL2s7T3oOI2DAGnU0lLqM4g1c0KQpuERXqSkZvwwsURBR5MdwVY8iadtLF0
7NCN5fjNzywKnyg38PgpBqa247mp2hbQLy+Kvnn4q1QOiC5haI+h6nlYrXi10H1ap6tZ3jFRoCqT
DNhVoMDYY287VwJKNu8AZfTx2w6PrWuZRC22yN3XTwIaolMWimuCxqbzLCQH8d2zxPKsd/U4eHnx
IhrW+0Ce18h3vS84VUvXhHLMTLPQ+01l0w02ScyNvUojb5sGCmI+V+6bkZaq30cqVOjZeldC6e2r
Ru1MsDyWO6sscLy50pdG7Z5XV2bag4sL7f4i9dCLY7m2JYbSsZawtYkXkXM6q+Wf5xYl6bQRM/cR
DClppJKSjW4GspxtRkmUk0OtmW1EnBG8qx4SOHLX76K/28H2rhY8zrys1I4Wuz466QJPIJiiRU67
ZhNa6wTiN8dajYczJ8+lv4DT+BqiJgS8ahJMVnLc+tmjXUK4aX70fhuoA1PKMnzJwDbz7lRZnexB
YhhbVgKnsvm9opelVs7G+m9E1/kXQVNkYrAlf+Kur/ONPkMNUdWUmV/bOTrzVgDgTfSn10J1Dk1t
WuKYcw2fmKIR6ZrMIHVOURTMmdMWalupvm6YxWoMcGO7eT2Ac90s3folA0zLe9g5hzMm97E6Sqxo
uuWv1ukURdMtgCktAHlyrwRh+lnUOcTYN7ODxRU5fgxqc02CM5H0W8t6EeypkbeSi1vZ48Liv+et
rvOO9Jwum/P+PqjECaVciOYwGkqdLAy0SqVWluaYWbUzGoneTY2OGzsQZoF36tlM58PZH3N2PWn+
dLHZBupTlbd7bcs61WorYNom2exjRhxxRf1VzR4bkEl7aSruX/WO1q7Xr9xQIdG+lFQVC2BINYlk
HeCHtMtWgQ9XiJklTJEzSnWY4q5NHqDWF6qPc792RIH+wT8N58fRKxiQKfk1JK5fYJK9CiaFSIqf
kTNBgJgzhxKlnXxrKfpcL9ehu+E0HAfjxxLRPxNWbzU7QzzPX6q4IfFa3utmPbwbjMbqqZePmLb0
dfkbp2o25bjZSTsQ2FAOHHBFLtlrJis1GSVixvxNr1T978qrBBkydE+9RGlwADyuR6Oyt5suY64R
6/uKxEUorspwNl7kTzvjFRHrjGFFv58v//dYg1kNPcjFV1/sm/X+8A3LWlEP+ti6q/Y69bTnwy83
KQrOeEI3LUeYCoTiRliobJaEU5CU2E65ryKhfERqz/IsJaCAfcLSpmohVHQ91K5BAsmDxrb+qjy2
t0dKpDqhMKsfbYtuyzpWxOV+ghIFcICzVVsSOA2hSX08RmVGmRIcMXaBBXuA82So6vxgtztiH1to
jkFss/mF+hoQ0krM8iBDHpiKOCiq3gjYWaq5Jo31SRC9213c32qAOiuqtD+xchA/SZD0kbPERxlw
3zRkBjLf4Tl6HaeSLVjcMlg+HteAz0zNLngSrn/Qa7yUpBF7CWPSGh+wFQsuFltL1Lq8kMeRGF0a
3VpZWBv0qUxfu7d/60x0FdQPJRtLc6/2MF71QJ/mi7vo6wnFfw4J4w/YaTaf81yU+HJRv/0r/LQX
rvwpXQg5y9OI6jt4e4NAsQu/oST6XOLYF9s6K+KGgFzRWUj7hAjcpE+PYnyXHTl+mwlFDn8VHYmO
n6REFmnLUruZvOIakzL+yf4zfgxMXjONCE3CxM9uSF5Kbh/06hB5fEfCszTK3K+i3em7LPWfYVea
Q/Vm+RTPiKpolPitAwkvowb21ZJqjL9kQoDDSRAzWsclZxmhlbqJdiGDorxvZQlx5kCJJ8v0FK9H
cBskknecXtwuh8g20LxkDmNfG1tJ3EsyURXJ0OSvaCOxPhp7oMLcG8zp8rAD/yZG5B3717Pqh6As
kvKkNZiQDnFFcNy17eEvOKSKqQPI1TP+B9hGJ6L5K6PEgTFU6zvNsZEqJ+UnL0Afc47vJd1N890W
XQnUibq41R3uQIPF6mqN/NZLbSyi2Jy6nxtuKpDNntn5P0IKK5iyogcmaIiznXl52drQcV40foUC
OI9uqTEx62HucwYWrNbvteHehXXmxHUPh/l041fF7BjBqkk7rWrQ7ZPrgkCHef1O9owgkQjHWxZ4
DRvZKn8ETOFS59jTHpInrfODLD2FQhU9ahPy7AwUD0PKmiH2QfaGnlbwXNmTKKqcdkQOrH7YlrpB
zKPu08yjGGKuA8SnsNjlxD+bQf8OVT3mxK7BQqL+aPaDaUJy3mvZ833o86xC11eH5DLYl6cdmPXV
hhQllMR6DGsTd6+R/ucrkuJsTv8mSg4QnPQ4H+XLZoFt6triO5CuIQdf0RhekS2mEwm64OO6hGtS
OdubHQQ0MRDjCO630NJNbspHtFrHPj8ikne9rrAhCvFGaoR8gLTikUwJHzOZY5E22v3LiCpusLLG
38DB9rELbyw5xmpFpFq6rYv8mWgk+IFWSaPpo7+22+18zGjcTZgIosoA5gJf9IGQyovZiOu2qHLY
paQGQN1a+b5i5cRi23SBGtbeoeG1ZGXNJhYKFQmfMtZRExwcorJGrHG4GQuU07Hsi1JID2W57xrg
bFB3oWWiYPTkZ8xJps18j7/0xOeGxYTD32onbxiyjTeKNMieVR/hWJgaUNQDOwm1dBq5LHn0XL0D
GApn4cgQZrRw5TGIlfxFsjkbpqLrYI1JfvyF79aXpzO1olXivIGNVZ2Nv10Uu0VIsVa8Te56tDIF
jgdhfPejZQiTCO9OV3leJbVCx7JUthPZV4bBRhAsk7T7lR3l+MRY4eH9p18QhHIi59kD0ezC5g26
Pu5T3t4DhDruV1KXOHc5dtMCtdCMIRsLTSu0LXBQeubT39976qK910ngsIDPNYVT1bE/eSwAFQMX
5MAYo+TOp2t0QGvBNAvveX0lU0m0WADQ0vuCb+wrRDHltyuxvVvF/zJODDOpaOQKZto8YIB3Z7i/
/L0tdkVTAXVbj5CfHuUMJB85i16YN4cGJpZ8npwBfAKZX66/hTjSgrbeWTkrD3WU/2NAfbKoitxT
3qPK09L+0Buw9j6dwMnfqdrPga6VRKt9pld5FWc5fE2JIJ+nRD1xsU1VatDv7KbR2LVfpxufBpd6
Xu/aM0sTT0xxZLB9hVrNOuCz1FTA0veYNbn+d5iFJqKZYAKga7TOZiYhUXOFePaSgfHCaQ5aVIXT
cOsH4Zur6FILPHwFPqr0JhIhYfM6H0uJjGcWOR8EOq3/v8pxWg2zSIj4gJnvnLO5+sW6HD9HPnkh
aWqGQ5ZzvuMoYNmU+Gv07Y7gHY0DvdwvRJ6fv2fvnBWozW6tRnTlKVRcDVZmErv+uYfDk+CPLd6Z
liuBDzQ2cpNUrX+MFWQkyceadnnZkkyZ+gH00X0+zI2WkL1uAcmEQ2/ExM+LB5HlEHsTSttq6VzE
7Z/NjnkQlhrHR0v1ZKL3rzaNjhTYHOdfiGjGkpc/zajVrSuYPIiRFOxlE8TiraqiDfPguc2KrBXN
aJAKQbOo8voxWt5WBDcyhIHsMfG+RNNOFVzeF8UP4f8TGlLHyKi4yZkz2PvlezIn2weK/qgXq5PW
ZnddfsFLOXCnuJv436Vnp1kxdE35IqsDD/xbyLYnbIQV49B/sFZMPcqMlPiXuQR+EI1Oob1fmWJ+
yIxzuz3/XZJI9qxSPUB3OovJKL1MFhO3bKjQqwAPF17pP1cAOmnC0iClA4o7kfwA69mDb8wHaSu/
jIWeOYMO1pe2DFDYNyINBA0AqUdF/kNfzRuAi2xMvABl6J5HY4ImR9z4U1ZdV/dQOcspU1ZItzXN
btD7LuDwvBo/H7EhT+KzjmftLhkYJTTWj5I0kzP38rQJtBuBBT4fg8i3j94R+hYqs1yAOSh2DEcY
hoNagFkxRnoRI3VvGuuEBcyGD/vwgZPRNUPgC5DIaeJ/8zVOVncI1zu5ZjbP2xD05Ae6FD/RJIcp
d2O7desMYt7+1sVuzWLuuWqdHXVC566zjbbYkYvU/mFCXh/RjZ1dE/cYBW32Yh4V2Avoj505U44u
/UffWKRygTznM4HZggdmnZOEUC81UokgCzECJHjdNo1qEGhRWct7cDrRJHvKSFe2/XilYOZEzTcM
x49gxW5btLTQDCoSRI7nf0DZs71+dDext1Coo29aqqKjMLneEt9F8szpMY2g309sNafKtgwvClY8
1w3cPyW46xS35KSX00hePR0BmuLtrie/GW0pAG6BDTfj3PrGyYptFzLcUYd7Xd9qxCAQaPBrCKKh
S6kWlCzp8X+/+gPkjxxkVXmQhqP2syV/pkYlXDa2+axES/gfkvVMVUFssf8yMyyCaWa6HDD4i+ZX
QmfUll6oTH5MwOUQVyAnQEv21Pe5s4DWXDCwX8ThJTgih3qCb2p6YJgnIpouIKweUAg95XRaespG
DI5gndeFHtKJt/avaVh3Irhjq6yEyeAUDZwVCO5lQlgGC/kriYBrZuS/poun/Q4FQ1nIG3p3UFgv
DhdCue+xTfo+GpKTz87WuYLoDHAP7O4669pUhOYWVJUh9nNdtKs30dYGNvhz6/sCJEf5eRrkNSgB
Ex2DMbC8PtSpWrkhCo6fCBuxcRJkuUKFPDF58Y9bMmTyQuBsUBobWHFkIkI+xDMVsqe1730qMOox
dcEiz50Pdk+aTeDhalvGHWqbRc5YjNRPxQ+4+IjmhtXQ3SdamP1JatcbbtvWwsDaSXFf/1D0mTML
sXs9zShKF0fmpcTkmN3uoTTwitpXXULGQpmUVPfX4Z4uxf537TKdM04GswEKOpMlP6MzpsDXAe8k
abdcW4uBF0n4BKKFHIQoy0NOp09xCbVIkeEWpe8xCAGZuXNp3M9gzWIY64HWTqGN5zjPG0D/j1WP
4QDUjmHVSLJKY1xLGaJCWCkfj00teWG4rNuV+IHWPXENV59TXKFY+FLZSBo/TeyxMeEj7gObZTu/
UNx1DAwLqs0GqxFpghyZ5yctc/Q+2TT/a0SkHt7BsPSmlKkOqC+fSzliFAZ0uLae1dPYVO7/p63M
bMpqQtjdHJGXXg6f5NfHehZL0ZyF8hCVJq6voZzNYGcn4UjVBRlpRK3WDqtDLDIluFzSIh1Izc/8
pLrzrWXyhXkr2bZablkew+ZFQ0mCa8X5N6dYAOhhgSNVocIWwQ9VV2WanKbPXXxA+zj5AecpOCWB
oVNVJ2FPaIJf5fqokB7BgCwzYbDJK6K02OR8Yszu1fSj1ivlr0uknCms2cq/xnwAhDiSAxaPKhAQ
yKe/slU7kpsG68oxxPiUXioMs/tOvQJHhsBHaPDLnhR/ngY7cR4V/6W/9O0++98+ARaFK17ZhHE5
Xe8++EbKfx7KRml4atvBxl/3klbQDy+PjuFyrdx6utI8FFMgj+AwN02qIluFFO90B9Xh7odIu9A6
y8BMqGN1pSoOerftyBLnPwJ7rcIUXbsvPlwsdcz/PKHsCcQFPlcsEPIfF6YO+GyKZeKti9w0ZQ+E
+0ToPsWdm1o6FguaslI8JyEITcPYlZE0+Xxbdq/YiEl134Bft7RaI6GaDtrrbZBGyhI69bl8x/o1
D6VE7xXqAxcWp7YjtYX9t66zNoHW95toxmsMZbNI8pqq5AzjmRZ37qTXPCTp9ge0i1F9as6Nuk27
RRImR9YGlXWoW3t3DJM3+WhWSO52lV+ksAqdXsfJLyTrYlKyD+LAKJQ0j5TK2N4MGEViTh6yuey7
19lh1N9/OzkOu1VaXN1VI52ONQXU1tOtVDsblV7eidFqDvwo8lwtW9yxPCOJblfxjzDgW3s9ly0u
XnpO+Pw0GvGM8xBtVmPltRC03gE18y3btVmMCB/+YR0i689b1mDJbpKG40QrqBeQXVCC5y3WUTse
6qmN+jCj3fpnHe9GNlkGKul1BRNDwtHVzAgUDhEI5piWpsrFs2G/LrtGDHn4Le2gCn/lItINnOHI
uCniznVinxcT1PGn6d2P1WqUv2W3m2e7XZd2SqsO62AeghA0W1A0Yf+lC4SpEjte7arH6YHiLzmj
tNQ/th6djgpSz3Wc78yS8oF9rfOclMvxrgv/Q/az7vQ3L0L6XA82XUszZrJBwkCi4uQxSLtdKX3b
0IKuYiQgEFV5rkcmqhjryTT7kRkHvegtJyJXlgaWBQ/wIUwJcSnSnS51lcr+nJ5UC50UUpMxLk/L
9pU0HKlhQqoaFf2P0/tZ6m9ptvY45223uOd7mNr8IHblltSp6jPe/3Wdnid9b708mdTe7I7m1Q94
78QIrCDpXxW8T65pA21Oz0g1QIwVnfMUsWwdEKyP7/kDBj/+vB2GDMGv2n2xlIwDDj8aV18NpKjd
UsSLyVVGG0zWmr5QFWdOHiFDeO9/YGKbyM+0yxzrLhKoHrGhmw6/9Fu5q8vUnGlxSxPJNY0zDXJy
wqRkPmfcJTWnsTE5ODMf/AhzKZsx36pOrq6mjKumz+qmXAIyJMtMUYPVHZ6shVCeEu26oPYiFc7S
iYUdaMSTd0qYJa80m3GDM4Kdf5XKOAH2iuINcqHIs5bey59wm8SZojgHTQSDSU8IVmviChXOc/vh
pbiLq/NWxPQ5QfES2GODl9Jnn3WAL1rYfgsnW0NrAhoLg6QlQ59wR8aDv2ipHi3aWU2WUZAbOnUW
nNqpP3n5eczozXncxfz+FCBlgrQpAYDJUmLSIi43E8OU23rU9bIU0ZHfCVk4SsWylYcqGTIQJDb9
QM8py1OGIJRQJpV14b+6bD7yfB1sTQDfiSO/71QJqTmrJRG/ztWcLHkuaPJtSBWE9bwUOnHOdiXk
EjBxJ/cs3VgJlx2iOy1O9x5Ht0+Ns2f7kojaKksqYDF9PgxvSl56j5hKpJZB+sjUguwjer+qtgYL
NG8xMfirsWuyjgKu8KfDsFS4Z6iJXQPYCyvluk24LuDZwLN0WjH5rGDqFupgqF65KX+59puNNDDx
eKU4HIWHG8aD9BekWkbyyt5PS3Hw7DMGh7RafhMCjq6kI4/VG2/zPZ+/+e6MjaEMGlr8rj4OiGdj
igSvFKPmUnrX7FhJFK2J7JfYaT1NxeBN/9nPs43ftRD4umXdWNjlRrkhwFr21u12NTbYyc0x5ZOk
NZnyrhoY7Cv3TTDNEhS1d7z3QmHW6APMwvzJwr7TGYnadacwyQeAtTaByYaSYPQEYFGL4Y2blp89
jxLBkjER2J80jOOpjB45FgLjYkRyGP00gFJl2kCNvyq3DmAeac0D0H1SydUXXFhqaZNSL373LL5P
G/ZM2RIo6ZZFtxfmOTpckFENBO+LJmOZ2qcUXfEOwdAX0Hhdw9oH8/M13m4n4a6QFElKFVhU+uJX
MwNYQTsDdt2JzGOQZ/gbIaXGR0JZx4N3K3lETdHqIpucULCUdAaujIPcWgARAdsINJqHkHuZMkBY
PgstY6AYrTyZ5dgGFZS04gCYzon2JNrExHUSKS8JCl5ZfPHQ6BZMA6h0MVLsrXeVt5Yc+xdNkZ+3
qahCIcJxoYBnNbmgGu6hoZiLcxeYpHO8FaLvK/LWAMWeYVgnon5laDcGeYFKbLrzKF+goZAZ3mix
/imf23xifzPwdC6K1Pd7EvhUcLOEShXTvUi/CchFCKuiLQSwzDQEk/lgjrb8kGjArTfnGMDvb+zf
xb735uoLUYNMbwBL1lhjQhDtQUurl915zKqLerbmr2xs4a5XFr0Eskv14TRTUOF6/WmdZ5FqhUnZ
4gHkDjhfisQBwrIaVO9UDG+grdlKRRCTa/2Vd6WcENXSfwv9vSubCAxgT4M2o5aPpEgOcCNS5Psg
nZxxLyF8K4QMnA1avGYN6TemudVS4V9l3QetNn3DivP5/xYbOcH+7QF9as+A29nbAUVXFWJppNzl
WngWfnRkhTqts56hFbWEmrRJS6wS0RTxUmn+n+t1+4kdkyJGdRP2baNrmFSZCrJ+OEaaWsBqsZJV
gcdMqSdN63FurjyjO1M52zLmLXVdwACB8nRzSae7RvP7p3GGvgi2Hm7xTLt94+lHCm+GD9i/OLWB
gzmcV/byJXoaNLV8MYFGtQC3CYwc89ZYAGD9aM0+CUF4/GhK7JFu56dunpmdPbdjQKA/mYW8Op0a
+vYVy6CnZ7yXLqPA2nI+Zv9DmjW8/OXNSN3H7pG8qqRrCnYqHM+K7OKE2WeLrRJUIItD8Syh8aqc
wUAnayfQ7H2sZlU8LncNhOKKWziULStiO0iqdze+A9M5yMAHudzYK+IqehvTCwfzkw30SmH+fxd2
5/UjDUHce46Z13iVKxYsA2E0TBq6b2/FYLFFIhEmYwTatbgPCi81Cu7vMSrzOVXZm/1u+eWhJ1Xe
1qCPogVeUiYpPDzpz9Hvj8xysbEh8hvLkqW/rPE6WgfZKx1wJAXLIS/HmbNGcWJ/HZ1k+mSQ7xQL
ChHJQ0VtuFxX3a17isw+MPltbIHHVWgd/7UIJR1zkOWtvkKkGM1wxskEqVdUnav5NPaezXrkMP0G
qu3B8eLK8ciHf1BREi6SGK6QZ6q81v7NuaR1IT/mJXEe5h/J1ZQKPrOW1LPU+Df9yrBhtX9ypQ+3
ILgFiKL2ySEu/EaWlZ9cnovSoZBD28LSoAO5E3Pl3hmFDrWcCWvmuf5wePqDNF37JNyYBhSzpY5d
6xFTVPW89RJLbTc/HvvrlVb7NozB6Z3l2G4avnHqhYLBgb3wCFZ1clbgxRc0RYcBNMV5OY8FohiV
8vDzrUtOtWAqSQDRQcftPrPa4wBBx0i2WBhqkiJG7tnIfQBgd2vliwv29cR5AaNhmcsc5sLM56O+
YYL16niW3BJxj6iGbnBA3N451/vgR06mj6rcTKjTH+WN08sfDT9iv+oKbaoti+lLaLCefom9JCNw
yTLVAMVY6rGFJ5a8tr41B7xTXyb8cnA8ZigjrNWJGygo8ED/nZHrrkiZi/aA3//Qi7ohreF0CnnE
NUHDuP2vK8KT12KT5Fx+uiy3It3taZUmQj9uO2L3anfJFJTUqjccBmavzYqv5kLTIt22FLPgF/rW
3qasKQkx3QwPlOWedNun31KiGiInFUqW3MYWRsHFE4keolEhBnFIC7uPM7C9bMiw9JY04GFISsVc
UaHU8kvcwdiAtHtDIj3F0cTBomms8vA69HhepdVpCDblnn3RLt8z/GPr4GyTrXRm5YWht+A26U3H
DMg555dQ5YyVNE6OGOUdFr3dt/TdFD/G3+vrptf+0fcq7Lj+wudvhhKpd5+moEb3EZljA0QGc4R3
cwwezrYJJxoei7A6GYtHXixDjTP2EfsuDzvD+MnK6CDB1KIW1Nc4P3Xzo/PnFblxPBwMnu1rrfNV
PjWKr98s2oB7BMwP4KIn8KLoeuGmUqpnJxNDiUmXUXmiEsJaJe/gYeIMFSlNMKkbwJc/dJMhxTEx
JQqQY82pmCVtucpMtm+nSEDpq3PNp0IcrcIFtDOIG2+PMSXRzqcd1zfeyQ1D7aZ+gsW58dPgBIt9
5nKM2BaTh0VeBTcc44H8hM5cq59U6+TJqP3/rf1koFcH4/1HxUYw7lG6Ml1CIl0LsaFipPOBGw3l
VyhJoRivbsO0scV2H1KYMjCOAKY6oOEIbV1ePYZ4bnH7MHxWje3CkCnyLeC3zx0PGI5Vm5+mdpzg
U1ItqXeATFCvPd52J2FtftB+tbBaq1ga3vGz+oDp1wXVW6Rq5xK2DDZ3cFP4JAelHLaenBatMohX
pdcUjFncTFp6kw0izvDm5GF6pXxWG+i3cQYSRM9IV8OoUNwtSJ4PXnDbLX5Uw9uBKgn4mHrpd9ox
t32s0+zqUgp6aQC6XJ/ejcFHQs3BrTrjVyU9ZOAniGTyx3e+2ttXGm1ga+uuZplkXz7tF1zH+MqA
O7DbE0HopCxPheCI9M636CF44NvgfzeyjB+ZzXW3GPCbsZ/4KYPB0DQm72CgsuMT1QCWsM9KgG/3
3kDgYkj/Go/HJP6EzdhQP3QV9OZOqa+Pu+xW8f51lhUIceVpX+JO/XxkKNVYZF04aZ7nt2KrCyMI
UCc9/34bwEZHEvQQZGKC3v5aOkZmC9lk56eHp1/5EX7HQGkgw9qj6qgd+IbF1T9lZFApAGEG3R2L
qaVy4lLDE4CqQGBDTNezdgD9pUPC/g17bVmq5SZmIjwYAEb0vwzf+Od8+upG1hsKWnIkvX90Xcj+
KTpxvhPbVch26sUTsgneEnwsKOp7CHHS5VIxoTcRVgNx3ofsGYIsK0psM9/mIMZEWCaIaAXZCnGh
mVNlzg7Rlc3DVwu94POvwEDLZekiS4oqQqw+W3m0lHA1qQioYLkHwru4yvPvM66chJrTwe1dfmAI
yEJC14N4ClGfTzHXGSQl4vVBg4EfcxSRicDkIhvO97HRI4MpDLfllW41MHgyCYj9ZnYnvm6fqTiL
EKDLtCxgBfS++971fLphoT7IO9XazUDSj6fNj2MjqEgv3cSAdJn1I10ToLIf+ux+msWIMrYBqtXs
xjFO3LKDw9manS/CYzkMKScAbUXE5YoQ5z0Imd4GQUAJMTX4oxNmVk6y+DVwyImcB7FsArs0XLhb
hxyoA0LcWYB/GQDSEySeBPuYcb327/AAhV8r3gccLn5Jt5WGaAr2p/sWecVDRdpzp8ciaNvJaSoc
ToS6lKvVKcrbOVv0lOSxBE3pcZujxYt739SyKykZE6KYsRfPhT2s1NAweB1ivNo0QK0cAgElZGBn
RlRB9k+b61E2KJ5L0rjVNqMuL5Mefj2wmbkKCi147oyoRDJm+yY6CF7s3EvvBrWmh917uIMLQZmr
KCzhCLXJbuCSMsPbYpd1F/AIPkulRVw5EeNhyA6JVoaZU7BOFy7tfP3TN5h75IYVO1K+hwdcpp5M
mzY0oEHsuduKlreWhUSifJ4EtqjIfnIjZs856KV5SGUtdpVD9mABHpaGbaZq3JZej/ll1kEZGVSv
o4LbfUmhkSIdKF+OnfHcIoQ4sBSVNwISE//K/h6YEwpMPbdVtVhXBEncqhQBHoBK7DdvZ+U6rH5l
5D3mmEo08PPPJ+4/+2HPZ1qboql2ofi5DwLjR//zobDk+ZB5/cpGx1nS22t1Iiz20XhxOJNJMvh4
QRi5f9lCQWOrfuyYbE2d2qGbriOTCAUxuhVNvjD6tXwIHDvssb6VvMQmfsI4Q12Q7PsfNVbI6IYb
LgHSzuOVOZms2P05d8cbUM8j/55vxSIMELdLcO+NpfvLaXaBxNVwBTKIKwkC/CYYTO1rCijOSx1X
z2W+QeewpQDK8RDn/ghx/NGLE+TFM5IuXPP2vsQ8WbyBX4wLoEcYxCTuBx2RM+u6OUMb8sJqUA1k
ivAyT4ITi+tGqLKcUPFjEhHdpSYY42A5X7QfEw+M6ZanDD3zZv96vy69y2gRK7mOBZDkJh3Gl81l
v2mqHv2W4Nj/MnSHfNNl16XA1gyFjbY/cxSJUwOaiuuJKJX7WEj+gvvC505AbgRax3Luz1VJxfNR
JZ7ozMhzyrXn1ih1WtJ9mFCXY1JJdPUMqCB336fi2Mm9uG/e83dNDpSSAukpqTVNDDIMqvbaRESy
FLLKkojRGPtSfIL39qHkII4TYrOdnMjCH/CoScUhQNkD9o0MYxKw3ONY0VOSjbzOqQvF9iAMfa4k
2+3J8NmHE5buDjDl7G5nXSQoQ6g2FRil/3HyQNIkLsFq6Z0F6aVkt6a9za8JvK+FjHU0lwuz1bgx
g64nZiOSgrCfClzpi92u437f1sugocY5BXBIw3B/ysrHCO9I6dOtccHRecwPYPFzlTBjpiKmf3sG
BfeyXUax1FtIquCcTOPmVRoDcMED1F8c2aAIl99O07J55T33W9qsIxnzueQ+iKB12SBqwsPGaZFV
xnYZClGHhAk7U/Fz3BKPVALoP5vopB21++SI8mtaiNKx8+BEoAOyrwGow61g3JIcC6v/yKK8hhTY
8V42OltYXHOhpyy/yoj0zrXyOiYaDSESHVEPbIU3Lf1JIE/kDB+a0L6Fjrldn3GEvqckQwVbf3X9
awCBuOlY5OfCk7mtZH9drWu5OamvYK2DjBCC1YmIzxWJg9+WgozvzWlU5D/C/JjtFAFpD/AaBuqQ
7rXcTlbZPXNs6YsAHiQzKmG6X1/VdCeVOCGjvaeE21TsbE/VgzAvCG/wQI79bGpXc/KujkkoluuE
rWig/2z/cm5cTkMLPtsOdvI7w16RRSAQkbfoGvibXciBw+RpKh9ja7BSwDDaxV3x3AWFHWrIxK4M
RTersAXv1DlVqtSqipO/4TG12an0a7rW53q4HE58PYEUsTkioVYJMXjosyV52179bVBA1dK92mB1
424whjDQmAk/PZ2O0UvekqZdJo2r8K1TTbOXW1oGStx2Iu3QL8sGOBN+iQalbhMBAP85lhLPTUpp
VQ5Z9GCToqrGHMjQ6drWzsBqHMLLegQqUuFatijbI4PSx8dKRShnYZOwIRhZFsZ0Q84qVAhN5jzr
loz0jOCM5Va/qmxhJcieM+FVu38WXTpIqMZ1sosp5+Lvi4DZTu0WQG+nlo25WoRZHHTerVUTtQOd
mmUkwCwZU+RWr7qOqoSgh3b5ak/FhkONKZVMSL4l32Sy+ZzwzmTaqAzgGSUvac8FKqNwzk2Sbqc0
TH9qUzQ0bvUldb7nI9TH835DQwHsOYlS9w33viH2IRv4o9kzjYnKMh7bhpvDLp7NUWlJ57KseieW
L8zoyGCtViN4n0/fVpqazvCIMkuNBqCfi8QII/0yNRkbghV37wRFx4aB5Y0x+VAv+m8Y2gVpXP8m
z84M8vCr0piOCGjcJ5DvSBokdGgCuV5IaJan251at3B0SbYixhgX8hd0u1UnHB3L+COG9wP4IOmc
3aqEX8nntE5bocFLwSAcucELFJ9zQz3kiqTnbZA11ijuWw9+tdqVoSuk1TJd1hcV4g7p8CpLRc/8
Mg+sLzdJqffsix8/CkMvZlRTuesbCqnPa1tvf+AhY/7AcAmJTZ+i6uL5CfOCM9CyyaYhTS9AZESQ
RMAthkg/J5w30SXLDVYCdwAMxVeGBsqkG0cWqx5BwXKkjX7ioeBpHLB02ZjbUCaPN7at1F95EWbr
IGMp1sZqAWbzuReR8W8oGJVA7vVzzN5ra5LPbYZU1TRX7FM34Y/HZTeRA9lXcyaTVGQPh8zBQSjZ
XwtHZCumkb11r/vrG5XrOeEbLRpnawyqcjv04vvylMM/ZD80C2ZddHXza5pWV1sTpn1UNvVXkCaC
4mNkN0omR76CzyCTmqXkvbz6Xurdu0nVyngJewraKTWsjVL1s9CNfmyAXTwZJNLmWN84kwYadGFu
pOnXijVHYp1m0V2BPP7XBpwfS3cniXBZIxcuAfyvGrh88kXHwmo67+Iiov9WZZu6x5ekVHTB9gqa
/Ax41QXBhnBi35+Hpw1DkCVyDsabFeQV5wfkb2JDqIcfLrmhqXH92Aeu83RHx8JzdmIK0IWJ+5OI
fcFk+h3EGPnwR7QjpOYLqvJHNFl/GTQapmJLVGZwR3C9mboL8/CaL0JAFePVPoo9cHL81jJOuIqg
S4FUe1ZCK/t4TWS6HaKoUF5Jq3kgf+nMsV8FOZPqDqR655hIangLM6AAQzDlWGGRqNdWH5BXGxbw
4mr6kTxrSW+yCUP+J0YAdb/n2g3q6Id27Fsq4RAkZ6BQFMNMKsLOLKTghq3tqrSfjsrfmMX8yBjf
ALYyqYtjGMkLEdSYMkFswBBMwLZGpc1xOVJMOOlnsmg7c68GZCBGUd+hwQtwlb6hvqoCRa4e2oUu
EvBElhLaolCZm4T33C0OJ9WSl/sayXuQgCxprqohUJHNZW/jo1qZCHYRJAahK6ventyAQtlpo6PF
mRBNPHz7bkaTIDie/xwmwTlgIVIa+DDsiluSnVWR0toESzS5LPHm1JaSRe/X27LS7Z5SjxLuIzA=
`pragma protect end_protected
