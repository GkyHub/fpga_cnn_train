`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
KUba/82/Wuqe90wyuU20+pyrwWGV6jKdT66Hx2yr0JOr4yH0gq6UMcWPTqeCt4LA4/FGnasUt9A7
4n/A1OPc3A==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
RxKc/CXfWtdKc4JyxK+SVjUyWKh1H0Vi9JBKpj8gEWCxPjvyjiEMXLirGT9B0ouwgD/i8B/H7EKX
FS6UmyPQck3/v6hMjybUK0k71+VDWY0N1tWVeN0xN3AzP6fKKgxe0WB8QDpEvCCuQYmfsBFq7eRt
K9t4Pexj1m/eA667PiA=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RFbbWYBtmcgmhVgy22jf41KagzLbVJVdWPO0wRLCguVgz8tEBve560TyOT0WvLrPQoef7UQArVhq
Cyq4k7UMu6GzEDJDNzIfJEHf41xZd34fe5nRs5PJrUdpd/lc7WHIzBy8l03xxkOAV9NmqFK2YTo3
Hfegy9w7o6jAqDdknNvxC+XPjEbsiK1S1tMFZ/IXW1emvfOauU62YKn6KEqb4ktl/DecZH+IgFIu
Y+pY1QSdlUnbfcKsSxusZ+odEgWAiC8fz3cWP6V1sesp/ydAXnC+Cx7gpCVkQuKEtWaYEZvftqC/
hmqZ7tycJdmj14g5W5aHLQiJO9SXfa+6d2SSog==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OlHzjj8dxVLYTPHIMukQFNnKfEQMwtEIgXtc7VJv2AY+SO43P/u9yECq0T9K3iEEmBd3937frIR4
bnas8ALCs27D6JKn7koyGE2f3kiABT9W3GmKhJD7C8XgO4tt8SgS/6yiCUnFvCCYzveX99qUNVIQ
pwC1y4akmitz1MqIhEXklfMRp9OuybK4f4m/5FDz4vQZvsaUgwKuMD2AsyLxJVI0hxBirDpDNXnx
V+AAX+dTylTaWNNnbFCoVlezVtyRhI32EhBoS/cF3DAKZTDefAVBGN+XiqaJSRlAj12iyLR0ATWC
bVAaYT9oTwwHaAAJ9cz1Cb6a4gDRi0PzBqHdXw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
c7HqHm38CZq+iz75/7d0a6JtFJ6oGyfB4ANR4jkLyn8eyOTiDt3utkdvyGKFAPKMeh6dQUOlqx5A
Hy4tluUm98ahFDcC/4CAYGBP3MHbJJqpb/xOaamHOeqzWS3ofIu0U8kq4W3ZrpV8vGHpB+/7M/eZ
FO6eDlJI6UHCOWrJtp8QT4QEvta32d8soGNokmzkomX7pnQiQZi2XjuhUAAsniIlUg/veAysYrcy
MzpM9ibLvq8G/60vwKTvg3DZ1TYOZDzOWPoq2YO+H9ENRb4C9/QT64/gjUlH0yVNfX8NYw4411hA
sc4QrSIHNnLwrKmqAZWjvKCBg0oJVLsBSKO4Ow==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ISZzH/1zFHgeqeakjnzf6qb9vl1duVlyyDrOghIX8f6bg6Q6iM+m3+BlDYwR2iLTT4d1iHvU8j4o
U3CSaOv9fBYKpmIn0Hv54yFHQrLRHoT+3rNHYu/POgf2er+A7LDy+vsGakb/WPwEbEzSwnW1OsuO
tiOHG0mGU7WZHhrPTxw=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
XP7kSMER+9xMZkP/vmn7CR0wrGEvGfRWZ6IoPmhU1kkMgcz+SQRC8pHn+xFX8eRdZ0+1cOmN1lDg
pQWaVl7pl132BdJEOl/bniRx6jaHG9MYlJrS0eBiPNZPkdcrUiuMR6842LhCOLhi5xsmI1bMPvjV
drvyx8QvJgsIYm/4New/CUazP4Ibxm+HkC4NchB+wxb1L0X0tZLAO2tuuVNJ8VhdvJiE2JXcBRVu
5kFDghslus+1Pgss4nNTQ+HVzDf2YBLyEE3ZW2K1GFtUBmAUHgkF/8IZX9DrNSUZAY8J0xN0VI/o
it27nUvUkt286A1MhuPABg/XkQc5uSftG+G1Vg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135936)
`pragma protect data_block
SfcEmqcvJE9VXfyKFXpDynzuP1a8mDAcgPA1Imowyrtg3LC1M6bzHM3fwfDdMUdhrXSXChyWXF9N
9U5dxPVdE1txI2EDgikNroXHtz2ZWgFpR2lY2BWcU34gS3VKKoBKhIVzdkp3dzTfITRquCeyi41x
MprsLnKTrtApE6wqmy3Mm7/3a4hICjEqovKnUP8/TjSaEdhrrwoUVNwC0VIt85GL2RI0PPeDiCHi
gk0wD5jbwy0JzKXCoMCLW7o4bY2ZXgXFk9XKV9bAv9sQ+y/D1G0Cru+YnK8uSgsk7hYaReLOejB4
wZozJWacYT1TPrKtuP2da2OyzUJEfYXyyt549c3O6Ex5eCgXjeImEWcOCOHDN8ni4W1ZBOQzGMYz
yTGxNpEt53Nd77YLigERMpXVlAKcDGVdOo9GjsdAwU4ZLT6pWmLzRZGsVmPvY/S/a6r3IJ+RARg9
3WHlvkNkk7mpzeoDqK92jeBMvu6qrB1XShhbbHOD6b6gxwi1H6TiMjElxgQ02431uqtziXc7optm
IrqNJBICl/y0JNTxwJl37TCCWPcWXkVX4igJ9dpIZ1Kq7w6kvCIDnSQT0ViWC2lmILpNj40NZDoz
arcFLX6OlVt/UP5x8E0wPx4TkJNR823yK6yOIs1YPtiBTfsHMd6BsQFzpK8b2jFSQABqbfzK/G6w
zhNxA8gdfwSO/vK7Nu9X7mnF+u/j9l42Eo2/nOpNNjPoXay2vxgwnFrru/l1nNDH0RqlnwHZsA9x
gFNTdNklzkyy8eWv0CaU7pbCy3RHaH9jHM6ZE1ZGRPMteSIpezXD7bkIKNE8MpslzH6xy86bnx30
VD+3w4suLqoOUHPYOeIzziYrrJp+9Pv4pqmvYbkjWCDoTfjLrxjvXgVm4QYYBRpWWiQkwEtXjs0l
ocCykLZ+t+zDlgJFb8/OaY3OvjYHmppWGT9hNlaGN31mcKYqNRJK9HImSMEdyFaKzdZgBUDX1zK0
jQW0jz7z+UssH03Uuj03PhV31vyS1h64iQ+0Nh9uBV/tAjgv1kVBsSvHiXEP7rLkmgN1rC6t2TIi
ihPLxmEAK8SZ0Wu29R5lDD5qdvPo9P8xPKqU9WQguu+rxklkxomYVGdWMNzaiauYq0zqvQpG2eIB
9ZeRqH6vQ51cqKpKcS6kzZLUX7+NnJ10WUWnrjfLc/S47qamygoZai0yM5ZNLSH24xM1B8R3W1hu
xLpP86h2HjfhzQeqWsoh0DqEkPub10mJNN4o4vBQrH3EjqzxaCY9R7SudCfx+IV+1t5dxvmbv/q1
wps7hStncfhuQGjVwGqzDpDFtUsEwugGIflxDG/6DCfRQAxe0+93+xUXKjNIwIPPMcdaOjqeA1R9
2F/xCVLRgcn3yvNvkVKie35Yz/0vD3ZzjC7OMS/KNai2f168HaZzjclSZNNbAPQ6ymQtYpvTxXx8
hozpGdrOnu2q4quMeh2ho8/Dvhi3pfG9/xuhZI0ui18NKS1KUnkqAuc4FbTnYIJXt8An9AF+DXTU
NgQ2Q3pwJdrgsxfzOZv7RyNXLsjKTgqrl8EASismr7Oz6rnX/R55uqNrar1JBjOTgDMGxqRnPV5x
ONs6FW9Um5hvMxDNI0N/FSmKSLxYozf2lxD9Zib1345Ix341cKKv80OhGK4JLIJCkeEyb8LQsEhI
CeKH9A/Esgpi0rKTLyZ/1ZGibfaa7zgOwFIYlVuXTtyQRw2RLDpi8iXz9QGsr6cpJjSdOZqdiYsr
F0M3ifhPWUvtiJZ9tPEsFr/hH2jM2pNJ5vMXWi1TVgy2/dIFdl1oQdjqNdvsjunH6T/qjxQT4Zxb
FOOznp8w5wkl/Nb/jx1rJOi4THZVh2dWPaE9CDYV1eOnxfALXkpv5hJ07WhoSGeUrGAZ5WrAslPT
b/2EOyC88xKDpGx+HgosOMy0mEx2ds2M0zBKzyz3I41raewA7JmNZG5eRZoLV4+1SvakbHRzu0l6
Mb6ZSWWSG/VaVttHl1hZc7TM8rPPuUvil/GKIPf7x7bdZlJXkewBP0WVdW7ST3qY/MCWh3Hn9rAz
efkoiGJJ9tahMXVGnrUURxp6bqUQpkGVQl9OYeXrL6fgMAZTocknJZqmEvVeNlA7t8Mul49Dp+qo
8rlpW02BGweljnqVxzManZzPjF0wsi/5+VMm5fkWma+NiOz7qbvn9QTiLP1BMe2Aame7M0taIjAp
wk7FlT6Na83eWSkNe/iM/hVn+0U6/hDS3NUfxgAKXI9P7jm8e3NZB0JDUNkfTpo1YqkDeZmNyic/
kmtUvG1FAVI51flfJYZZnYkYGgFIzELH2nXF7WYqIOJEmzsbpZRcKFwjC6gQkTcgHjtF+m/1AB23
qXF8FoTqecijaYz3KK6m7GXScICQ0IpWLrtFmbIjHiWxYReXv6BJaULr4u5uC1NhEuBbyIOSuKwe
L2O0cKvHZ7/kcsp87HtpUXA4qGrr3e+8Cy36z9J8TUGV1FS348z7xG2O0EMMXUSDSzOlGgMci3EP
Sym/1OIW5efHeBuMZ9mIfBZJN7zetveEvX9fSHV6cbsAE1DGZesIuO7wkiHWr4hDWabQ3yMLAxUz
iljRldtdvmXM0XPdbGpnShr7RQsXgTWDv14jlVPoUzjGeDSZTOAX4FbzQjnk6SlSCSkS8jnSsDnV
ylkpUiU4mEFplQrVBiir/fvO2Xvo2Nr3WrO+tjtyLHA44oyS64d3T+V6iebXaU8AoEZ812RWJQzk
ChyH4tgmm9Eo2MoqnmobGJWB3/SE+PbdFzJEaqr0HwtYmNT/dwdjyAIhkRmh9hdRiR1RgXxb0tYd
UIeiDe74uNBcyCb3oB/YCYuphsdg9JIuwPliapNRDa4qULc3Y7tRUpJV5m1Ui2CgtDZj1tojlgTS
F+2hzNM31AqrrRoUHj3ihRWPqtrKMRK/4RKl6dwuF9n7yMIPmr7VIaBkBHCKIs3tuTUz4FGFy7jR
i441SBsnPX7gZ9n2Z/DapkYGmLTWoafIuM/H2F1GJyvaG7sNqgfSScuDZMmJD9QuQpireVIcxBh0
sZlMfHryRhG9/wg2BciMxZvgs2qolQx3WVOcvltmenVvXspNgh/pS7UUJQTZwgCOODr0blmi4Rm9
el52HgFdlsYXZ1W+y3A3WGrTQ+fr20EidE3PKCqzuOawbj6Ig1NeIViq2Oo6VEq8cYEXWLdtOjbJ
V+qQwiMbFCmgDaNL2lr/rtM3+Vi5RsXtVTF6gzh3snBYrOvyT4sfaPpxWPLZKT+wL+F0P5HcLMVW
CMC89UTtDwDlvGW1/pohqhdpc8U0v+qQ3I8gGjfNfHTtMa5zKg67ObJnfWMHE9EaJPY9WbZrKmfY
5wscfaFcfP0t1vh106ULYB6JKQ28izq/EWiwpGY1cv8tC1SyP77/XKKrRmxtuuJqgp/Z2uSsygFc
zfwRuv4+Kn06dZV7aCK36rk1C3jfsjYeYGnyc/dvQ2ObR2b+5Cfcwxl9fYBSvIhdfEnKS6gO7xHQ
InOrOTozv/vB0mCKJjLN0DrVYKBeiNaEjpvEuQxKhAxqJYAZ50h4ny+2QNvtqrqHF/Qa03KBeu/a
iCZGnEaYbO5XRKAR4lL8s5OVay0QNs5GsniFNTauNNT9mCKGrSwlXpngZafm5SowfCwHJTRa56ic
UalAwqZAbAXZXRAKjE2VQWxNIi8vwiLz16MYrWY0cXhCBa+SYLZT2KF7fFfM1V1k8cPtpTW4ivGw
a+mFwf9PiwyH6Gg18XJb+4b0YIavMRHp89oY+rrNCmFw4mYLe0U2pBjr7OLTEgAbDp+ofl+QlDWv
c5PnXuXA8g4Un5ZAuivFsgdUqYQm/PZvCufmEWVZAbU6ZKQdLOLpMwydQoDVPtvnZCUmKci79ZvN
FNDZN1k6oh76FrlRXZetj5Lr8re+HPuYpRyFnW+5bFlAS5KocXefYNbWyhWnBVCri1tqukbKDG1W
cxBLOUNiOvqe2ibUnqTzC63KrpjAmbKYf2v0fb4b4UBsM/aWzjcg2J0p/VjnEDnV2PXBTGjcZAxL
FSHkomVqe8Ej1m7h5pocj47vvktN9pAjb2fuxeT8pGgSkAIeOAy9BKci70AxBbWKmsHbHcbsp2ED
wejaKtq05SvsmDJEyqeeSoR3fP+PFOa68xiUE19hSp2knxM4CZzQEjDmEXl8kzcIoOtQTtzMpdOv
St4zkhxXnxOWRUcSjgEqReZP+hgCvrsQb9iuJFjYzv5Gw0Dh3DjhkR/he1lk+XMGIgyxcK4Lc087
73OCxFl5YVX8BlpplgjKSWofdWNKELComh9gEiRkfBraJ9QWMLpzPRz/oZvzHtHG7cUZrYcpeuWm
5yrdup3p6QIB5bnVPgQctvvVcuJb5xveRgTkJWHV2qqH8DYkN6joE6D/kGmYQZxf+JO6EjMbRMxK
S4Lk8PWFcBD9Uoa/l/rELletcRLdfgEYJOrzgA+RtiqA6zHNbvXfiNQQDg6zaC9ki/JyVo+Y3tZi
YB1sesOmJUGHDf5NyrMgaBWYcm/5dDpFm0igbbSdD9Khg4MXKRH3EyGAgfzMuJUidreewMF9tGAv
s8B9fgzl7P3diM/TsTkoMVlGqGL1EjGMUKGUT4D3bYglyvgHjaZejrhEJREgoUX0ASj+w4siXD0O
5MPF/Ye53Zu0sZZlxyRIVidmd2HbKYy7dVaalNNvLQOiUpBCp1pyf4XjWcFG71TWkUzb2aPFVtky
iUIS4zR0z4p20G3NxoEftgFy6WEgh9SMIVoVMyL8G/CAhR5xzAlZQrbgN9im1gKH9FsexB44c9Tt
XZ63zlj/QWwEde/NjaS5D+WvkBg+kCWSSsKN2mdGhPbbMlpVz3OIq7hs66kr7UkZbSutJ6WpWJnD
nJTZV0fdXzAAOxwTgnULKcxqX6VtUoM6fxngiGCngwsxT6WfxUtRWRXurNBo3Q9iKytCLvaoapaQ
YJpRw7zezkeOJUXgsYajBDQTsOtZs8YAV1+R/UE9yYzyTPTDuiBxpoWN9N8dE6mzR29MSbi4O4Jd
xKUuAuKgBeXrR/rZjKDdvn9ww/1NPhRr+oqiqA6HccF9QG4vVRcH7Z1OtxUoaz6Fd60EwQL05jkG
gRdlMH713qAfkfKxIl8bXLIW/X4Gb15XzvDhMIiauuyYzmsElf47bi9T7LPvbupyRH7UGojsTHCh
fM7YTD1HZ1hVc0/SYc7fw3S7k8KBwlmyD8c9bXqZOkEJP6/qiHydJEY1zhTgsMcfedp1sXIOd59X
Rb2tJfWpulfZbIL5QHMlv2Z1IWlxT1BobvcEmp4QKR0nQkbZwYkG/GcC4z4upVKcFerVZw4XpFr4
B1IBstYkjN10VzDH0D80HmcrOQwMazrpdoc5TyP5mYF9ebeHmsKVK/Ap9y5Ato2yJgO2t3eAEQOt
ThpCCE4R8WOQmPsdPviaDlAofcsVwQACI9fzZQTO38Mo3PYm2LBP5C3UmOlH6S/GC3T4mpynISlS
UzerJKZAnpanVZCj/eEGfmXxg3vB0GheyTV2H3SJNLUMO/GvjzN8vF3K3ebN2sfF2mosenvfE8XA
0SeDgA3nqjHP2nH5hFOFCNzvtljTfq8KvakhEH1ELKOafsMLdxnM8q8ISL4jseHqSifMUCt4H0vO
PFxUhZU0NoB1Nwo9oJpG2CZEpsq3e+mFxDZDFcaUP7MeLYoXgOHRyMMOXuYrMJ9lI/3yQThPoHdT
r3x3P2SKbdNtWy5dAjNKR/7mvSaXBvjIDe0pWitqejOD9aeV2HlH7/iBMNFaIlddv54lr6nm4eks
vu9Y7/JAoawNxx/db1t7+4BXXzFcuNpmm+dzkE+Ugz5k26uJNVzvfdXHC598zLGTtVw91xxZeCDu
Xbe96z/wq4KxPcfQU5wGPrRYKr54n353z3/UgxWBmBMWKhrG8wpIpGpK6Q4dK1dfsc8K1zhTFcE4
JrSELzo5cKR5cMj9M1Dtgee/5a0nLLGG/cKFLZzejeg5jI6lrwfk9w5r7nwMTMVMRfb7QBQ4O8rV
0DgVde8I1MV9cm57IKlWHRXmMayMzqnu9v8ohz9WVp4vy7vTyyviFeDGAX2FlCovR7nNWfOksnbU
zsbfn4MDKR1xwnoXjHacGplkVMhGXRJGb8jDzq+XYZZM+5Gk6X8zJzPu3ck3eYnwBgeWyLXZq8sY
OAxCPRbOGCqvurAz2lt8fb51CbRYF1DTlAIfdkxdomxq7pm1jZt5FZU+y1aAvmCzdmt4Xqe0bWDq
/XNZ0nbqKGkOcWgy73F4MveatQy6E2Bcdd1EHLfFSCGVE2yEjxZQwGRQSSykePECCchdILHM8rlI
8Dbpn2OzKiMEr/0L3WDyTemNhJ+0h5pXsjV2AIeuZuhx6aZbhsIRkewzXTbllp0eAS7Brhtirt9f
/W4Iz3u/svtcyZiy+VYUYTqmuGI7KLIMqLVDeLrQMSb2sNh3OnT/kBUdci2GXlcrq3yxw7vvsx6I
OzpxvrRnHKy84jOh1wo/rt4yxbSyyBR3ePFW2JBHkRsoa+ygHYBEiBet7G0LvOrt79DQHP98zbiQ
JYRSU4JJHC363JzMrjUJmcOKsF3rnaorQAXqwpp1sIvvt2MRMd7D4Uh2oFtU/5K4M6D7rw1DU2+f
GWdtwyeBaqju3GDvDbqXr8aILXqk6WcD9pNkteulr92Ys8na89b0Avma07SITlQc6/z8QNC9e+W1
Rzy4cLQXEBbD02ht8m7jRAXjsPY1+ECVA0yFNfHVBujUK77kBcsX20S2yxu1mK3ToqeNPPw9ROhf
vy2+zhJD9ZRX2oENudsUGTz0UB/m7diikaX3v8mjg85oaXmbTqAej+siD0mAENmsVzBMRYiYCd8X
v8LhpQlsnvaSq5hCWDpvUuEjmxdsi2VPTuoTJ3SLJI2tFQXGVMxNAiMtafEgSt3jedouwCP6kg5W
xdC6MlRMUyNO9Ap8VerDwR+k6drwyXleEn6ZC+A8amfpOyPw9V1RtecH0jx710W57jDLwxRM5ky+
cDMqu3UZXvJGjTzZmUgLIn6uYh/r/UbmLR2u5A4akNNTIccGKy5yWogoIClLQXujMjJw9TdMs6sj
XmM9f3Uh8MiFdDYOjvcG1+WQJ5kDoL8Iy1pgBqCF1k/igsLMHkAtjvgNvLFNFP+3ONRi42ZcOVVO
JTSpjiswbE0mOilgwFebvmURAuFPszntxNoJaz8jG3Q4EMQKKpMQbgYeH8S/5sFlGmge2sjMgu7r
y2KhUpYZJ2Ew8ZTPs2ZwJwgcFmdCXid8Tfhhwzvv0d2HsY4TsUrNNjzgNNYtH4N6j7zcTClFAndi
XIjR0wTLP5aTSiK50DVVuq2vXS5la9K+eFn0xT4mIUbdJ21rgGpC67fdRyPdUhLYQ2bBbRmC84Mg
ETl5es3SuZ1Mf4K9jlwaXIb3lb/A4OA5sijArjlfATiKFAGeG4DQMyOowrgYF0+lpQi933xkgK5E
PuVIt3F5pkS3U4BZfutcFKftgaAXmSIC4vsuAoGrW6bukQB1BvH7XjITaznyQ8O/SvHkRMMezO5N
NgXWpOeSkfU1M0++BrZS3Ix/wtBLClNCApuIzCHFFdpBYTM2b8PQHDNJtQIttSVUX/Q1x1ZAd03j
M5wiwftlcM/kFXfQ20IAKhM2PmL57kU/3zy5tHvAcC9QiXu102RhPwvkf37IXOoSZwwkCz6QJyJI
0YspWu3x87KeMBXKCOw2bpXl7j30R+9nPCGpXr6dyrcGrjCRZjhalr97qyGy4ogQPYlECg6qiDmV
zk/Btl03Kj/69MHPtmy/iZBTDUeue6q8MMwohwIltcpuvwQOWGROt1LJ3dGrE7sE4oLfF23Uwsc4
aMtP661BhwKnH4z9gDXa5mav0xIEsfXcQq9PvBjZyYL5M60UF0U/DNgan30yNqRvmRoTsG4te4Y9
5LHbDkb1uoHC59/2Iety1Pp3Bb4FIhcgFgEmrP65gk/8a1k/3cxblVWWlV4h5eR7zF7OK5XXBnDL
r0zCCjkT+bE9/PdKGewMQBtD8qLoFlsfuOm/0WDGO2/hegCT839x5gH9mHgnTSIXKR1o/f2Ad90l
4DKp7+3ulsWELAeuPna3cZpBRRCsQ80Pz4e5rdw0Nf51yYXT/U2T8lLSS2IprOsDV+CC162SIkck
UFKagld7DzlZCHH15piVrgzMBU1+Rs8hagPicByKyPyfMZQCnVuxXQWzgqdGkHfwid893YBKx9oR
2KfQKySzosnEa+1M9cnRifKdmmHubmzifAUs6HnHLjMB+jIGkC2VuDC8za7irlEeEyPWBP/D5gC+
OtJ0CBjz9pV8x1UpMc4PVPBomQog65OShHhgiVXn6f2lrlu7kyxFO4ulp943M+q2UVemWO0DbnuK
NCo0gxIv8fYnn/u44tSqZ3QAT3+/qlZL0oNZRJjbruCrkeZxPIcqkJShhObBMfDKHTlW2+80l8PF
Os8Ap/hGL0ypiWCUu9iRaa0k4Zde+Osz/Pw3dLlsc6BiIpjpT5LHZt4ACo+U7N+TROgonbsKV4tO
n0Pu6QtgatJ1iTYoIcWyRX044xb7JSyXlpbkDxrDu0B8RPd5wVOXjV6PKrb1kiDH2PBS/xcAu4YX
z5E1SqK7rkBgcnqQbifM1hiN1XrUkbtNVhzmBA6KmPBa3yqspsTfwBRjg0I0lQ3jWB4+szEiHnnx
gFpQmS2dcHJsOO93kcq8EOYbCvWnqVj41znmUGqS+zUsROonf8qKb+ZsPeUlS20ok+42ddi6AU/J
WnY6+6R/PCKjw5N9a3a8m+FdvDuNWJWQTJ5ghnOpdfoUFrijl8vbJaRKMIws2fzgYTZzM9hDE3E4
CF04Y3fRetDRiZmifAxIls02sOEIwt6HJYDUSVIMsFCEixddhJ3X9GUTibdp1mpmOl4KokXtxCCe
ZsQWbkLM4M6Pr4ew/FFRPc7BA81mH/8nk7zsTZWEIS/Mg9LuHVP/6GC3hRdGdEa4KeS5UQAVze7o
ey+DZMuGCjayS0MKTE7eTWowYl/DBFKVBaiDGz95v6V/LMThVuZjOVi7PlaZpesdpmN9l55TmFx9
HotF8iiu3pia4MJ5rixn05Pi1X3tuxv5xcPhISnfPTRZcc0o87BsbD5T7YLfgSFiCVnvlqYl+3iN
CbYw5oxIiI/PS6D+jPnqGhck3WmbEPH5VZJhMz5uj6FYtrKxZVffriU7JolvdhzatSqITPGfZOpv
3K8IVoDZlKS1Zog1NA4VgFdmF40F3+KsK9SKuacGAXl+V80at6xqEtozn3QQRVan4nitS1nIx5Nr
dQgi+NI9UOx07w9xDxnRuh7k1x5AwsPX4hJgP/pStdLLSj6DFyV3pemee1z2OdYqUZbMcqtJaWrv
BWy5NKj/xjXlZzGf89wWMP6RXbuyxiLaKapQP8qxW/XtYgbcSIsbX5ZFYlAg1Zb/zNMwc0YvKde3
pcA6W2Pu3SpVQdhvocE33VbI9DFiMry6ECU7xAYUDIWxepHEvqfs2CGsZWEYlKgU+UEdZ0rpLCYv
kZsHMXzm2CPZf4Yx8VtBGyhkweEQn89hQe227LogxMMH2CoxzmEWPPYhj+WAE4zjyxaX2u6TF6u7
zc2xREiE6cwx4Cv6vMaBoa3P6wM45b4LKIIQc5M3h5/GZYje79alZ9ApYoK8FtLcN90K9a5qhHgM
m9Vqkz8hcCLWZg4y/nJUKeYTuv0UuWftKTt7tHuoa9V4Yb1ZMuW+2WLHHRRfTKDMrx6hdG3f/6yg
Dvpgl6qiLTCwFlWaLAuah73ogktJAGDMcCd7JMevavngmqnN0KiyN5fAc1QmDOsB6YVGeIu/eRze
3YQRR+A23RAPAsDMXfiCGDiaGEYQrK3QXH1Ibli4aNxHNOSAmJEER9PgMVK6Gfp1OKvvJZRPIBXm
IgO/tIy0GklJvHAngMQrsN13BGzCgXFiYf/Yl2x76scki4wVOAmCJjq63kVFg7t0RWTx6fVZeXjm
ixWaXS67R3bhr9sxGINWuSnLEnUuNcOwwbEBm7Evy2fCiVWxzkePKUthz65qSKgKe0GJLiBcFOE4
MwIavLi65BdWaA0Zd/QuSeycymyIwh8H0KEh1ljweGcOomw2XZkQriGQvRzZEHBWdQSLJHe5hIFe
L8BmvvUvdGur0vcMq0VsdXvAubaBNOb9otwB/Xi5BD4glcW95898ZWfS3O+IrsvJlQugw3NgJAV3
6YFlSZyhr35r+54zZ8YNgWGLmQyfEamibvP8RDA0yjl3+rWjY6NzXmpF3LC5zGc4MGjAzFgoYbUN
pT47c84g0FNDY3+c+VPuiZZpkK6Y77aXj+kEJ/xW6XZLpkOm4RLRxDcpFGpOsaq6CeTt4NM9fxyt
y7FsgblTnoetgxe5A0E74FV8qsk/3BvheMwCxT55UIGaT8huZeE+fosIz7OeOTctH/0Q8yrx+otr
3DFn7/J5U4x0KlIgbzbbndsqwyBkidNz9a6QhY5M2lYHqmFG1V+OfN/X+5EKgyFlXGDxOdvQ+/vd
yggJhyZG+yljw45kfn9OCHDCHk4ySx4rycrYJmA8KDMYG5tjj7JRqrPzJlFWxP9S5HOnls4KLboY
m3TRJAOU8SwuAqXRg0jwlyjGzg58TqIbadQBF+YnfYSCGhxC3jre28gmJ0y4X8wmslbKBNF8/gvO
eXcAK+We463WhmryDM/sKr/8X6nBmR+uaP5kVlz5pzBlfKRm65D8x5z/dQA4Ak8EkwoJrVxouKJv
H8/0PLA8KXWG3DfcMruIfVIFXWjNOOu+2N9xMVVwdsXlSNu4mGG8PDr5V5WbQ2XICREdD0UWCnaR
QhIOnsismdWyv7cia4DpQG2tFSNkGB9bpe9OH1IctYHQ0+r58nx/TO+V/35ctmaD6KLP55RoLirH
CiUs0eFH4ajQXu55b69h8ha1CPu+jvPbzKKxIOYmnrOs+FiWl7Ol9Bi8YnYbNf4hcRy7oQzBX874
Wbo6nyb+Grir6uh3paZ4szias/UlmrOppos3otw+bpACU811SH6xd+DZQW/Z4n5vLfVnBn3UvD3u
TbdKrYJflTs2GSe7rdSnYtoUatQm9s/dUCsLBYJILKYdtnYJreh/pYnUYhTi62TPXovp8jqzDKbw
+IPZ6TKSM3wBUigl0H7j0/mjF07lPOiIZcDVBlNTtVmg0fnkY1zcHZDcSZ6o1zMNAeWnnMw2cjEH
gqncIRpU72Bs64HjN5B4Cw+Slfs9g8M1Fy5VS1BT/40iXvQZoD900TMsX9fAH09aIwcovitFbK8d
K6Xubv6hEzQi95wp2i8ajsLGo7VtHGpTneh88wCCVjwK6WW5cQu5+bHLUbknkKal2FnbHoA0eXtG
DFCGUVkIo4vmtSCtPI72oioHDvNVnYWg931vrYn3UcsX27UfxP2ggEfotUhXMY/JpKykYH0s/VW/
hHojYVaPVsgktlxc36vlT79fFfp+fP+iuQsiKv4wWQzEV8bZoouWNtaqBxeT9o4lDYoijW97yWeD
pk5ogNJa1FdX09TDEHhg5BNs5Zrlq0MVni2cCi3Kb5R6tJADuYx/muLtaNVzn1XvN+sqsVxb1A1J
d7AWZUlM3xDFXGetmj5mAf9JpRS/syM6uDaxwK48unChqUdzwHcrpOo69FpfRwJCM4QPfC1AQ0R5
fZcjCuT5OZiobIkdyWMXrC8C85DXQuR10GIXtJHk/sKEEC8eVrSGIEym0MeW6BbBfobGx0gYEfj5
OwLyWhPUoEHqRFrgfRXjsmQvg2CwZIPpC8vJFRN2kDa3Bm5KCCp+6Uqlp6AFD2WHwtnp/CDGR1eg
ILxq0mr0fjAwDbmuomUg8kQSV2i/CKcvHk02Ip/bwQsAM7Nko4HM+LgKU4S9JlThjQrNgZ4NB9qC
+nQKy497Q8wrQ6sR7vdimhs8/VACkt8+ibBLUsd8pw5n3U92UDUcRnkuQxMhpVB8PtyDt3WcS2QZ
5FuJ+A4DvJbM6Mko9l5LgkSkz3b9tXXp/PxgCVNo0ajjVYtA1QM+mc/oVLXoOtZxKG2iOpWG0axH
t/OsUmlKC050RWerpnEzgZO9A2ugMdBuS0dgjohhM+fLYADbsm7n1fd+17C1TOYIjnxdr8yNNQLG
vStW3LpecYLIzAvPWBcJTd1UjjIoPCGdBSBzCmbC/iaXq52oQ4h6qRJ12ct+HoB6kBp/kvWCrrup
vu8/KUpV9YROc0W8XoEqjX9grf0StFu9DWQqo3OUzyH1mN7vyJWvbIwpf/ovfqyoSqkQs5MPPzWH
B2eVbWCrfMLYAczx9Yc+GXjWN9fKvT/fZU9eqH09Pq+rHGw7ZlvWHCUdTamGuIZ6nl61WSAGAKAQ
4yceVd6+tRxSGoF1mv72UgXn86WiADKXOhWzVcVNgsVcynaBWfVCm/nvBuivEG1AyA60n7h62cT3
sX5OuCBUB8abrwhsveF7yeKw0H40eK0WK4Tsg5C0TyQXZ7xkglisP70HEFadV/NjoD/UGe1zXD8l
6R4A3XSWUZRomWrJrGwgakPCB2z2bwgjdkNIriYwpwOmoa3LB39PbqEJ+g7IAA+2mX9qRjKF7Ybt
QWGxOrSvzDAynb9jeA71cdWKWATl6BWlqA5FsStesn5OZTbPPHf8GURt6v7v5Ny0Fkr3KTaf6neZ
4DliWXdx8cH5JrVA2thSGKYScLVlw0xmUs5IhGIClQEfSvz0pULR+GRTs9/RzsvmlNrB1uAT8lEp
I0QgGabp8G+u2UfXilbuYewnjEOLd1ORhXV2a51ePHI1ADL2pK2RLju3692SGshdOC3rirN2BR5d
zP08ogLDMefffs1ctNQJ3dlKWgVNrNNJB4cKk3yWIed2lyHYc9NlndXnY5uJaZ127Kp0Br8iTLxj
5Vo1bnDcHTzMrCREpGoMYj+kxXll5IACQF/nQP0806L3uD+/7epD+DiLIX6KQgYHwPDkWtnM4VB2
WpOxlPZQcqNolQ/gN50KzXTX8z3vVjwNsaMmZQ2gSmF1ApxS7CihSn/nLSkWvMJ/1E753P5ByM8g
PWVS0zXypkuiwxJTHmccxtZkF8T0Fw3gZy1XEDQkYQ+Jn0fnIYd2R7UqD3FBRea/lTpYAzHVU9i3
duJ4Lch6kZuGj0RK0VRr4ND0xmulytKak1XwwrrK2BTUKKRePFUWkdfuVD5V1nirIHjuz10rEM/A
WManjKnAjXlB9lZfFY9jFWSpxGXynNAh5reEkzZV/KuiDbzQ9OFeFgVon+1CsYjIKaYhvAE0rKGQ
E2ZcibqYdrSYA2SXB0YtAOTi1BfKNRQ/+cq7A9i+0kcqOfJ4P4MyCd6UAo8Sx1905KYIGaG8wEuQ
hZ1tbmxXsCeoUfuKrePuKnL/+X7o7LjCvdptCjv5Oo9hqgqDUB8vtJhJmIWY/lDNak/HLcR4PgUT
aRbvV4YQ1tqBEW45dUThRoz0wLqN68JncakMcEziGbewJkp4ZeDOB4HnhrptFFuFDONfAC9rh60U
K4+Ko4h7sStUmWt9uYYUVTPbUOdlLzotO4aTaEdPakV4tThDltgbOuWlalrI42Bnc4dA2SmXUwBE
j3BPpZzXQp+uu8DdYNy5Jli3ySLabtLVT1QhI9VVb1PN6eAYQv5OeSp9pgryZZRYF9MdBgn5X0EM
e3IcxTiMNTwgwql/czdhL3v9BAGI0y7VDC0pJiIPpxrfgiEG3WlBTQ5l32oFhXXH8GuvDc/+iigj
t6Lj6S3DZoiCn0Owoi1uu0et9ANr2/jxTaMia4+fO5FwqxCpyfr4RYnnJk9fH6xbttpIsBGyDJoI
OCd0pCBwm+Z+H2AoFtueb5zskLBRjRHnDMSGEEggzPvmDyFdWRIq6f0kgLBSsZo5alg5puPdiodX
z9NfgfZvt469srxAhyMR5/eKWVF9QP4jm65wnzY9Y8GRVGtwtuuao+CDZhKLNYY0duiXk8A4cwsg
LYw0hfslCs5aFL6ovaYQ4NVnry0vflRcLFjVLWAsgy0IHtiKYjFGMJvXFAuTmaSMKtqlKsYjJubV
OEhrfzOIZPhdUYPsgKru/dliGUY2QcHkwLN0w1OsQuupSZ8gwQd/WCHULhE1crOeIV85YuayPZEU
bpHsWu/U34w4F42Zft0J37LUWwph1lmOlPwOP56RYE+BUhZmaexTYYViNa+UrSkieTCEWoTt4EVP
cAZeEdM8ej7mBfqrEKsO0Rj2kNDryUujGxEdUIdPuncCE9fvd3E1M++DS6ok3MVWNwPTb0acHVSC
5dh/8R5J1QqpnbEVtn0ZT3Kt6xgTbP8ZAUu5aAGuM3UiuahGwR1fkJWIoSpUxvQZwy2Nt8Dzc1rG
hyGLrlpUbPLgRvBVqjXXj/UvPYYqZIJyWJHv8+wfoJXuoJKNA4N46ATspFviuDkNmWy0Ql0HfEa7
NMNVbtantDi9AMf17OWm/+gOjezQB5kAo850bwReqwMZuedRcD4OY2w3hXo2yApORyUb++NR8frB
81nYejKlR9OdgAiuWCsMJtotA6ClB1WF1iOfsJGpGl3NZBFmwiG3A+UQ06TZx9PahgxLtGCKbPNL
qufPsi5Lima/M0ycNZrKTRgr2QtRzOtK/iZXm1ZnBY0f15JP/cvhTHMhsYLRiD5fQjv+Wx1FVQs7
ZOxnUFZyV2vwExzVGe/e2UCuCEM/rzJ5d8eyQHnKtBbnanUETZm/PZOx7EGtys2fW7CS4E4Dt/Ym
3O6ol9fDciEqWfVc67O9+Mm7Y4xUFaadES2dVXU5xZ/92fgONSIPrAFwXxOR/UFRk2+jRrFMzE3l
dnv983/mV8PffCV11LOty9+hxa2336gEvlNYBRjQm1tivHyCj/K3C+dXA32Ri+fxEKVqojMHjfA/
RCLl81BFqV34CJmaQ0rluSStNiXjjFwaTnr3FIXx2J4cuTRgpGnVDF67G71a9GkP8TqvDQSYI6JB
Yue/Ou/zB7k3WPjlWY6p+/beHFIX9I9zcM37WbmzTywi7RGRBhh0yNbasU41SJYPd1BVL8gciMt2
e2P51ERhb2ikWbAgRYc8bayuwWzfWpg3fEE/VF/hyOE8N0wU2L9/ixlRh7dBniJ5FlqMJArGIEWi
3mAEHAsWHFrMmFXG5kC0IS/SFcgJM5W0/kkyv4/7rwVu5FnztQKrrlP7LbwfMGilr7WgEmClQPqA
0eVTztkgJVXayspdzNiHlYLaEVKA063fKDqkYP3mT/Q6qVAp+ORRWb88AZAAFUUEpzwmqWPmY6Qe
T1JZdEWjYuS1Za8aYIS4e9fIzyLFD3qb/o4MgF2FYslMmv3v2ouWXuc6FWxVscBSVsb4pY9DLoJ5
Fm/ZfXjiBW/AOufM60O8+goykAjzlx4O1bkNSUQxkkJA6uQlPX0MmXv5N/Qe4RTl3+vt6Xvf4HIg
eEaDnD7AO+7Jt2XVTnlpk/O2jyzeioe8NHy/F7f59OVkAjBbaoqDOjYuyMzX8JbcsdR99aCcFM/F
cODi62/+MFF6VYOsYEL50EM5WBcXxN+/S5o/O++Cs8YdP6yumlCemLxCYZc63usKFkfkpD2MAnCL
r5NXuVJ3w6tHRDC8EA2Qkq4ndaHPdsNS1QbQtJ9AJemiLULOK0Fnbf26FrXqYswPzyDokzXGbWN8
1gggNsU6p+c0LF8yQAR0FhPSyytIFoT1SsYY+SL0xrKqCxKCp6CVFK6rgHMviBsHBX9RtVU5GUaV
FMg/xtcGEK/cwj6Hz3HU4w9Izl7GdXkkpkOF1q+gDW9a9G8VceL/MGWhXl5NsQamOltbUq7SSzc/
hM7S+7VdVmSLhOv50AGQ5FBAtj+VPY7XXsuCXBRmuw51zpdpRihhbfyr8+DpZENmkT34BcZuhplA
aE8CuiLfGRzeV3WX2gwZSfuqkXThiuHt/yhwJn/Bqz0uRLEzTspQiAJGL3/OC/Brv6f+L3xcRWbA
QyhAzYjxjD3qcNlbXK74M7DeqmSKenZNxpgiGAf0OQ5K1NU0k4vWmaBMRrLl92vWSwwSd0ze/PPg
+rZltcMC6o5u5+QmW3HUaBiSMCUTkvnnNY5juyPLzH2irYKDY3Cs/O2dq2uAmcH9JPOicHbHGdDE
vIsFb2Cwh0xj9Wp6fzWIrusu2ShVnhaUS05U4QkuVj0ctGyR+7NS11lEmi4Knylv6dgtI7FpWltj
lVgjMlrQaEcFzFKwdmgQOBMjTfgbiwASx3Pc2BdEB6CVHasfwGMvr9V9U1bduey8dNbxmc8GC5IR
DO+FEoAW57vyC8twLasOSmF3CoqJwFt6YSuq8XAmiH5pZqK++ETbY3ZNDsNFEiPkPYxqVZFfyR+C
AHsZsgeDXCx1W6bBwc6ToVENdb3m5fz8SVSFaHhpb9O7De4Mrx9gMaVxbmguMGnfYyvOf1wKvYR8
g0RpeG2Xj+qfT74eQ3Pci62+dTvvQVarEk4/oFJNPthS7lt/xCjaViq39tAi4X0VdqbORg1KE0EJ
fAVWyntGb7lXnAGNZmj8xs4Iiu/FgMGsuXi1Kg7CyJJetp5TqJNg089oJjYqieWjFQIya07a7XrN
Rm8feuabNwDcHvBfQQR2fvmb4xC3vUZAuDJQDsM4wFTZYxemg0BGO8DzSKHjTxdImdRZnySrFdd6
f4EwSjr0cnV3xpyNnr19OEa+8rKH9DPUOmppj2o8r+eS8rcVJd9bhH1o7jUPH6jZwg7aJfrMEuCv
qK7d9kpLSDa98GIEhG/YyO4+nX/+RP/pAxrMKwWbGBc5WR23JzbgygeHLFTW6FmqKyy8nFfbpkF3
oDjvx/FevGOiI/11goODPL5RPmDyRqYi0MhykorZSw8jSRd5Q2W+SMSZvZdTn0qPFY4yJgZl1aTF
4tQp/MjuCFI7UDjYBj5wUSgpwJn3nlUgpBhqsYbFHGEuNhaBGtRHdjnimWyH3pJ41VDhh5uJ//nh
dwCMrD0BPILHDD2CjPHpdt1Kfz83uwdNFJUaCQ/dVyG8lwsFhtPHRaUsLxXW1/0VQx4Mwd9Xd7Xh
qWLBriP/+CEHyJ5BpGmIZXyuMfRBCoyGtRvGvpfAHMu2RwxojB6WVPx2uKdt8Ve41un1ReufbWde
h428Xb+FdglVrVz4u0z9xbq54X74Y3HnnCf1WfZbke62kL1il+i6wmdcE0xfLAf6s2G+Q+krzLlQ
pwwxxnMRiC+7PFTxodWPZIpJIg7cUNzmdxAi9gfrl/vpJrZxbi980LeQIWxTZLiCT+VvfvNB0o5n
oZBgqdwkB6IwEGR9dOExPehVfsGf6r1RvUtyHuCMdsSxY4ODfcPX1cgD25Ij/G8assQwF/uIWhaP
AapA4nkqIIWO0+sv3b7za3NUO8nl92dwYqMRA6jLhSj2fjoTelfi/jDRnt9epFqaIVUr1Eh5dVEJ
yLA5rYwAt266yw9f4K5dCg3B3y/M5UpQC0swcabTqcSVupoe+jisQKJvpH45J5sugqXdQMrrD45e
uKq5c8a2oRdawig+Jgn8VQIOQ78t3HclwvxNYXr+7Rg1qWgaeZ0DK59EJ5ohbnWHTkG9JXp/C8Gl
/9l1YuMWSDn4keWs/nIPTC2k/6tjYyg7aRsVJNaFtQS+D5QJJd8m7zb3dH7k8S4IHUr/k6OjiL8/
GfEPer16SJFLeiuCMagFMK21RCPm0wRuRieNzJIJEmgMsAGVc9x2wsb6yZn2rx/czAwGyGoSQVaR
OV8wXE4iYiTcBGMh01sSZhAOMpMavUatsFDWnTIorw/gvNG/lkvBiNu7cUaDLvNj5C/PwmvK6yXO
5+TwO60B2KvTnpV11NY7JdqzMP1fCMWyM+S6FROocUse2AZ6vbbmxiW7MI2AtvYkMlpFEOshs8+l
WW4vQ9h8W7DHbXhhYj5vsOKhC3BiJlmG3pRxf7i0juK08LXJyG1QJsDY87cxEa61O0amMsj79S8Y
1ZMjrEffc1RlVZya3Qzxdj40MB8O0HEOfwuBYfzgNhNGT5gs8mNjTMyIHiIPRhKdLhxkvcVQxOon
GAYDIbzEdxp0MryN2EmWRznhw0ihwpANIZ/pi64VS1yarg9stYPEXhNIVrWLc8poHyd9daSsmzHo
50W9KUTNFa/853smOn7XibHMwrJj0Lvyq7JrcpQd9neGuXR7kdG27HW/gYMYXkV87pR9VaVrZ0RL
OM/DHl4xLOhjBila4cbY+tkVwygvqMIgjFJRwwqrfUQb2cMRMd6ffLwgvN7C8slyiNNWTp3z0Fn1
YZAlDvYvFsB5Rr+jX4O/FjWPC1As96Mpot+g1W5OVCeR3uHPkZAuCy5a0068ewhR5OWMycB04vb6
4JIUAJK+pTQI9qpDKF1oBfqeReboYkrbXKqk2e0ZAtZvKmg0ALjzvEByZ6sZuuY5qeNByRn/S4qc
rf9v3yvc2g3EiE8/7htvj7oCGyyBhG+XTZc7odXCqYMN/W3XZI1T9jBmKcd9JOrleM3p5pGKFWE0
QGFICbcuLOcIieIvCTmeABhMSiU9DGsmWcGNC/WqsC1tRYEHy9YdTtqsylquuKPOHLLcWke+Sat8
+mn2NynWPrWTkRP1UBj3N3OgsZ3e+wsI5RVN1bfHY3jZBJivF2oSxH1zLFlv5W8ysmcjdIKUmDnH
w4tv7gKGKi5nUg8FbGee9PXo2sV2Qn2ScrFiNw4FbaP1GfNPOCGENEmetyeXE3HIeT8zgWmDqMIX
OFgD76eL3r8D0sh+8ehSPrTxwX3vvPllXCQyvj3uD43bCujK0NZEWrVFp0z8jaCvZeR4trvPi2hF
ee063CdKNkMAPNMyKPCU1LyS+9P7FFhtvSEWxBlF5mhb/f9MJuvpwjxtQNjsM7gkVNn5v5izez2S
TBGA8AuNPFiOktYtguFRDGkUeqUzs8ftP9QG4FNY+PzGVEvr+zbmf8iEnyCuRdxLDtDY+GJWeas/
mtHkuz2jlKbqs1IIUGqBI2mEQXD5rcYMIKdqNY+2Xta86Tobhy4LDe9fre9xEtOdbkAu2WllF8S/
3cq5xgWrnOx9x7KHvoGcQbNLNUF3XWWvKDn4zCkwR7XgDD6hOvyBaT7ONaZ6gnP+GHuJvHb1uows
hL8NAeq/I1kA7ON2dlWx7HIecptaRxVBfzMtaB+94f55cBU+zr4dY45m1EiQEySTul3MbU0V7Ved
FRctOwDNZWdNWwipuSphcLY4+LHC17z0srCNh5htgBHaOeTnSdGTH0Igw0AeRKJI3AZ7VxWNRpoR
oInRuwF6TU0mBU/QVTlwyZ8TpQ7p1SXQZfrGO0qSNKh0UCvEzCff+HSTh7wy7etX0tGB+3ZktZ2g
Drponywz3Ml20QHiADQsVD9R7Pgi4JyO/cIbQfpZvAHbPnAfXdQNLdq55B4OhOVHCbtSannxgFrD
4BXqisIYhbNbv3LMeThBrKt2HgwoIUwHwnmDOsp2dyd4keItN1aTTCDwWuxM8KIxiNCnGQfJpWqQ
VoPy2GwCpSw1LVYRQSvJyFxin/klYYzCu0pb6Ehu36yBrQMi4d2BjAc9Qa8TCDrOi7YqpKL5ioim
CqZ66uXEGlFmTftvJN/QyS/fBCYiTIQZUCkvdmRDThfCQNvCxnaaCH0VQAlAoHfYSF5CbdVx1xJI
JTKi6RkdNxirtGDydLIVv3BDDXJ2XK2EmxevkSSCrPzXn82ONszE3Ogf4txiM9HVKNJDrBhfeTgf
6CGZS/wktt6wS5bwsd0WAzSV4KoKwCUl6zBH7LtNq9zLl0qCT4mIe2w9tY/RuH348SjE8TeMg8N/
o/JQrzO5FxmFH+zMY3qfR2906sB/XQZZ/WrUZMIWdych9Sx3v33NG6lATZO5R0efOb47n3hGMJQJ
ruM+6v0ZBBVWpDPGFlbByBciSIqn4cCFedLpw2xJc8LAS6oy0woAQI6sNqCEjrcIvk6NlHwFWzBS
cNtoJ9LpyIHpGlNyKvMspCWc/yz8lUZnXdUvFJgR0uJpdHY6q88iVOPt9oSDmN/J4KL25S4dItVG
wrYyqgS2HqgyIwgCrkSKhbF1J8h7iSyZf/k/REKaUwIknD0cvpOKiw7AQbdRl6t0xh8Y9eilqOdd
Ic08hKwxhLKQJHO0TUpCY0yykkdwdWNXbRSvrrLEBO7QUbIat38ehGNo+Nh9fHJjh5rxunTxV1oU
AA20AfiZ0nVlfoyn8OIe1PTnAS+AcTtKGCn/pK5v//9zOtOHiJ5gOVMMNiCLzjMuwmrsiBze+per
+JSU806ee+GsU2imkCdeR63pwf9KdFHXwScqVjIT4jM+UDgH/7Dh2aMPk0HTGCQzrlILXmGGwkON
ln1XWGbZTwT7JN9t6HGxW2FozvauBn7YtAOOGt9yW3XoJLxElg0Y6LrGEnmncE3Hu91j643eIFyg
8oEHhJSIlque22xIj2H0jvMo5bJokITQvLSk/HbyIbSGkpZieuCoWd560AacWNW8xMnYNSUQMRF4
0OUPIKszAYOYutNtCLLM32P8wR00ShD11jzMZkAd00/z4GygneSb0xnzVUT4b4cxJfInqHvTGQkf
DXRv/urffDV6Xk50TqhzsOJe1OaKb5CKbgR0HN7CSDWo7MnDbdWm8eHhJg1fRWbHtwmq0pysDL8m
SetngmDLFqqxSUa0HwKc9t4/Y/B0Du7Y7p+e4BvBe85JjcmI/RnCby/PyiWi3ab9iyWbOGpkHHXl
HU+CJgPIEi+O/6jkG0EZyTH3F3zhlP/vODNFrSlXfdqkw/lbPR1EyuRaNIlgka3Jwugv8izmsTNr
IDFLHbYqG8F3slPr/+VNMXKtRj4GE1j88e3fAEF8J4reSf4Pr184g1lSB4p0vy0eJLfhUVCBVF2V
p406Jgec1hp/EMjpQCpxIBtwbZygYcGu48BCOtEeGgNlpjK0yi3zxbBMhX0x4IqhGqSzLFX3LUsl
5NQcTi858JXqC/6aOgzK19DI9hajJx32VZ9qH4GnyWs0BH7xJKmt99TJCULXBKL2n8VSOlJ69T/p
l1tLYJc9004nJ74ldkZ6ya7Nk8sQ0Nx8SjWv9x/e/Fz+FJoClr/eScTwxj24nlADdSpvGANFMt3w
YOnHp/xYkDUb5vDuE/ASv7eqlzDBOcTmvV6fecqTp+P1Qo6z8OrocBq5myTdxDUsC1uWeX14wa7f
CcyvIdddfnGrxNAqYdFClHv6ZudfExo436hpwk8Uy+TbFu7W9zKAd0dTay5EW9cHqWS3AH9PzLLz
7wZ8sfPGIFj2XmmWp/AFGqIT6sHQ1ZC+O2Q8IMsGKUznBu197p7mfKF0DtHfQzlHwDuPs9OwpOBH
3XulTIc3xvHZ6OjwCHhhm05TW6LxfeicGBoZ9Rb/ak28CX0nUD0dlNeUv2Db96H3yyPCaUGJThvF
Wvcnl9QuLTkWXq0GJM3lYnSDccROHY6gEoZscIYNl33KhvM0aypATDxDw6w4D6oiyVlQK3yD1yma
RcPbRe0P0O2aNY95cYeffN1Qj+Gm63qyr6qF0/eW5EB4HXfUFkF71imQp6KL/1nEDIw1KgJPaaA/
Iwu4Fgcw+TXX98uM6k/rs6AsuVbzoYLb9jQDWEQSLq2WO7mmzsd5YYz6GQUhQ5WZYlppEGtarKO2
E/TQJtzW3aYLPETp2HaNIum2b5AjlEYioxYKWxQHMtx+E7neN76hW1rB3mloMOSd4ibyJzN4+7P0
4XC9ZZ7BVAeyMrJ30+iG/RTiU43oVLv1PSMUWn9Pb9XEMXfjt/LmicplWpUjdFxgbNwnbf8iBEol
EASP6iv9OpLmj+jFS6H5ngW/pDRU2bvWmOmuxCD6foKK9ZCkmkt22y+E43DpmTtMnTPVXd6Rbd5O
7yo8rCBampUBILxlHn9E/AUxjZYKuxWzdAkyQiE4uodE8ip81M99R4399F3b/VH9l87xTkEdp1m5
JNs7CF4R3UffL5KpUpX5VPyP2aJwhy9MqpqcxqeWaM4mU3Ub63AvqhtQak9xkbPiwSVrcCmqsP76
fzZr75/TAwPoetW6osD2aXPyLfL+Ac++Fe/oa7IGqPlg8A7cZ0CeD/VOb8rUxRhVNgyhVHXsIGK+
B5PUW+LS0tKkwKB1y+BAEDw8uf5G99fmqOKA7UvE0Zyut8X36S3opL1pIF2JWgKET0otBrFfp6+R
EHfNdLF1nHxcQy8Chdovl5V1IeDn3Uwxf9GhBt9uDyecVGiTEmgw7COCgEtqGoR+gHMnqhh/VtYN
9aVpRrbpJRPIyIqnDIgHgpTGo4zoEEevBinb6pU+ngOk2ELYcvp4ArcgzPdRYSje3fck7Hk4B6Oj
v2TZfU4gq0LHOW38dmeCIRyK09FiB1+yhNE8g+3fzRGmj7QlK751TZJiPjdntmXKNxmX1A1ZfGi/
hpYECc21nEaN5qg5N54cNmblXsfc4XjN8AfxfUOOGqVxNQ1u1kO4dTjhavuym476g2yifY8tppC0
WV3EOBAEk319ZP7HL9a9FQCuIcucyx9zIHkJcdMRNELOrCdh8XKxby6sqCQ6kcwjoRAIkfUg3Nje
qWpaVL9Ssm6hI/Joo/3RtCZRxWMbpYV7oLz6u8jNq8O2xoBr4s63ZiAfJVdzD/oIpqlyoDxz688O
F4Iy70JqCTuWI9h8inwkEtIVDkJ7i+oxE4NUf6v0aKqeV2i1LF39Z0PbAIbq43ASgjxSxN0XRIKn
CyBrYfKhcwBXTppjv2Bgy/vqJ3jZsJR5PhiuN+u19WWOiXRft7wlDrRJ4BharW3elCvI8ExQsT/7
Y9pg7OKAqn4J8z+CeRcUDZvR042z15cWp8KRJT6gCfNQ/0E8bJn11VtJHA3dbJPBg479rUyFOeRs
m5BDcKpTWonINCRwJcXa8pSDtkhXraoWbGuSYdbJ5E5w7nYf3omnHiAK6nYjwjRzMh2jtzuHFdgc
mQAk2tjE5ThD46a5Q2G9A+xEYImRgFiB+N+/zSxPb0amNz0MtBKfEYg/rA+rgtPJ16cObBLH02f9
T+3dRh4FfMVcFQfxpIVt+6TQPqt2hkLTJ6iaFkmGCCTQAyX0RXmX6TXt74fJibhQVwU07CZfTkxU
gqAH4BHP+RWjJzNwzIoAYQkV+Ruh1ViFE4HeTzIoV4JZVdVlIsrZhUr9EOs1NhkR8jUU6bt/wnn5
K/tiUcfot8Zor5aL1Ao0FCsAEto1LCjqm4IQvX5MsEsjM65swZubFqpdoMeRmbGv8wtmdKQ6VvHg
PFRIpg75KYYqiSMnobvWSxnPf9OHJvywfEvAJ+Emr1ytRywJDXc1V8osbUTRZAgbiXY2a8URn9aN
0MlCaBam5211IMGggLuHMUh4EjrZV+7hn0sE15zKb6RoS4FWbxR4pENl8hfL+T25m4jANU0hG50N
XIfxO26tlyjO24y9f8FueHUc68ffJngqrTA/+p2pVE6mMVWXBRgB4zBd5IYRLvbJuRCtEAsHQahb
T9+UUMGqSANVQURqNFedGQcaq+WKIPUGi+pIv79xPoUApCWUgY9vGqyuTj85DlhyNf8vmlH9iEnI
4gVaWEvcswOxfEiUFVWmMIpxDPfv+Hbc6JUZf6+W0ZNdUuMjXZaj3fYABbnRRU7mkmMs6xDHpktj
jEjUQdWEmuHS7B6PnfZtdgAgad0CQvK5+S62uuWlzD4BfQQA8FpYr9Z8rE1CS5wMI5yX5m8m79hb
f4lUuuJb+B/0H3cn/aEIu4GmPRhbQWnYOeblBbniNdIbHqB+/WbufPPMKnVLSDsaikYSlVFRJlUC
Lg2Ff3F7zeoU/DxPmmgWmQCotBUjIGXad7H2+TVv0qWpGYJR2Ju+uWKZcKgQtMuTXG1hRhGlxH5w
vyLUNZm7foskxO5Zm+CjeU/Wf3vvSvQ/E+Eo5BapB+rRNuqHBkKMxrVbGeYnJpFkZESgeqKB5OZd
5X6D84KCK18MebZdeVZZNP/h7dasIZGYOPzuL0PwmU2DUhOn+vgloHlur8XA8OMiX1iOoAWlZsiq
zo5284cDyZaFh5guA3dqxXsKyc5gOjnFYIJ5A4eSsDCt+bVjrjEemTSutwYxARF5z4xH5juQc3dQ
qs1Mrf/ues86UQymJ6guElyF0n0iU0GxuxsgF935CRXr8lCyE+Y4YDJGbVYs9tCU0BRYhg+2CxCB
us6zSkZkNBiEk/1q4SaMtQdkmfc1eUegOy4xfK84qdmKh6lprqDPizXQ1JShP4VHOA7EMj9uX2eE
PrmEFg+Dee+2eS71bmKgghW9WF39u7uLk028pUiLQcT7DsVg7U938IjpLVlUD+R/7IqOesv4Bg4x
yQmQiKg6Zyr9CXlLU2IOsel1StFqojzDF5SFe0n6Gb4dkN3DGWdZvPw7rrTm5IJ+NVsefn9XMyW7
EwjvIrycLC4qo6kuuiKDQI2FRLV/pv87a4XpAQpf4rNGC7eVMBJ62Y7vGtxquiM1dT28/p65oj7y
jfyb5OsW+DHU3kL/qrLe/e3aI3NHOAsW8iBPe8MpaCtcanuZdFjdGzeSfj99iVlpaDtRG36qTjsR
0q0dDZ49W500QKTcCRHJoQ5Xg3QU8gPSLuvQKMlJWQtPbaaF2PF2bJGeSEC3VSYei5C/YJmEcES6
0EaXHn+9KhUbfATKrFIgrI03JTDTA+t3GOh1qz3pJK2ROwrStfmjLis61hpSR98jyI/GRD81uVtx
wsgPeO8Re9phawYZzxevgZ8RXg8YPXsSuVO8IlCWgU7q31K/xe3RZPt2mieaZjik3TRaMfWjXeIw
X73ryK/YXuybiZ70EUcASwoCOLy8lMbRJ5ZR7ylgISNkiqw/CqOfd1aFT6PB3BtuHcSWsI4lm3L8
nebjTJMuWn8W5C0EBQa2+jVupD9V7R7/Opg1+gwBZ/z5NKZjVBGNjhcE1bCJr53/IKsp6sklaAEw
nO5v2jXbq4tDge7G16JgkSzCzzNRAZCcizpr4n09CUSeNYMBmAAYcfveYirfXJxKZAjxWwkE3Mhy
NxFaqIsfo8qf6E1JLqU8T+kk2OAEuUEHn6p0tvzqTZBlINCsCTQwCkEx1BiWluzy6FJykPRZJY2z
I5V2kw8BHUAZSU4yH2wBgCgaRQdH8i6/W9UpzSc1sQxe9U5TyrW38cfG4vck6Q+mDrKOvCKMSn9B
oRm5SCH2R/RimaTdtNbbYQfoUxzuwbEkp/o6MKvLBxLLRHk/c2lQeXNHO0gp69DNoS7stBQoudHX
18w4aCj72IWw+lnYddgoFF/8S+KddEsDPLhCspERoHKRH1c9Plt9Re203a5AyplLbpWrqazj7z2N
n0MOLRftc/cqOOW73r7geglyVbclqlYd+rtk8rxaHW+wAlh0ULvKdbKg0dTC8IjX+P/4J9NpetEX
IQymjdiDpL66BMjiZVEg91bXloajlxUlwTpAlong50Yb1L8QyOghSBKCkeOE5pyd0lRJ7/rQMm9j
QEn2ZuLwKtv5gX6hsEeaqg/1Nlt9sZ4T2vZY5aPCpYYwnLdQJQrE4z/nTeJQUfYS0S/JjH2PmfFy
L7L3GVxI19DqRcokdtNJBsglhjRB2x7jJChh52A4NhdEGkF60NurQwQg+WWF3xHV3PnfAldJl8Ky
rqcxhlpE3wOVRni+BxePJUFeuCCvdyZ2txpCBiejDQ696NEuUwYbhz5XX6VUsamjNeXPAwTi+i9D
ES2jG+3QZsPN+yisjApj27lT0JIG0XMG4tiWlSAf+IUCzTuRycFspi0Oc60SkI5l2UbVT0shSWrp
OsTki1YsPktItBlmisbrFQ3vK8mOHpQRfsEf2NZG+hdcCGlHgY+f5Ac5vRJEi0nkdXEUEnWHcnkC
wCU4Wr4v1dWbh7n2vH0uFSrjQ+Wt7qY6ZEilJ9Hwult+QSNYbZeyEshiAhbgKmZGEjsf0zCYc5mC
/T594cgwLRrzclFkCWjm0Ze1SO2fL8qb2vSNK6FgUNEXZCoqKMliLCl7OaCl0CGpvs0NXFfAMpba
Jdu6JMb0qGPEwn59RcvMSpw4TBMLrG+MKzXOPVoV1eFVpRZJRVaeFFGpDCdCyN0kSEBfEpNCD0tD
rASC4UAifU3SzFg/9t4V8GvNlz9bdY25aDt9T3Hg/9jcLJycF9KVHLJEsQMi32LCV1T3ZGJx5s3b
vPQykWpJG1TMOccW5XMk4OOiuKbfi21o+Ejqj3aTyQCPiqGjpq03NyuhE+6RU3S01oh+nOHwoSA0
h787txARIe0dnYod09URqNL1dV0Ra4Adx3//7i+g8HWUYq1J4g/VIJYW8h/d0/SKVnvh6De0wye8
Thib8hhBoKxEy8mfEOpMm+0yxavGXpR4rFDjmBNmG/AUdHeA5qRU2TOjG+fGutQ1c/n/umMJ6itN
2RPH7LZfJQPAcraZUqOxsdasbFKrW0FRIfmUMeDWWmcB/60Q5q4QCecQiE6TLRUhTF5hXiuU2u5S
h6fhpb7M5fW1yMQVS7zgQDW5A1VETIAJd1JSRAfFpl2Jmeoq9Sya51EtxRAJpPdfPeoQ3x2qye+l
/qk60ZHsmhLGyWjxxfJkxGEI/XwUiPLPQzikZ2MSS961fUQqcHP71L2WbIuQ7mAjKCsqTgCY9lug
bzuvSfnZK0KJDcZi6cQR8QUajkQ4BMWTaLecDJLT5/ZAUDuDP8s7eJsEQn9pG69NvBfP6itQXmcp
d/PTqPpYoT+NsczeAiTvWnQnBPAPWiHsQnu5xgkaG3ngnicA8U2mNk+iC+oe8uw4tw3moUtdDafQ
L5Zf/SknKFgIXScbZnrO3XeoHKzgS2XZANPMfK5NMaI9DMehafmpd0k/IKrFoZhAH2jeVcJVFIft
slQS037lJ5CV42kM9tYm4x1pOpBpkHtvChZr0Mj5toPiwzXd6bAwWIW67loz6YTkT9g+AbClB5N2
/23wt6QecGFCVoMnP6LSO8GD8auXWiSJasnVAz4KnedeahwSKLDqWt6SmlF+RrhSjXO+C6xjOHER
3x/7bM1TaVLblroX3XEIvBMAIU//17pvpLw7ZrwaqOp40W9I2N9LRSfNCHNxgZJdX43t/zGHngID
bnQTSPyTaQSbvbOnhWm34/lXCea5CksLvvqCCjD5FNFy+hRbTwEl1/qWWeE9dxirqgSzc3jDCqkw
Velz1BLf3gBGjW1pdus743PRwP6E2PRRf5kVBcKIhpB4ylXSq1bsxfbsJZHGbqSYgpB/E9Gs5hwt
xySBg4cmBWiLdDOh0/Wf9kTYro8uOfdXxaXDxEffskj8bLP+0sR9jh2eH/TVaoYfv+t7dGqcrEBF
A0lPJ31cBs57iC76oaOQCQBYYmGviTtZcmI4F1n4HmsmJYI0sv+ajLVGhJ8RGMn0+MPoHqpy2qYK
c9Y/Jkd/ze7pcqLIX1TVKN+pn+kZkU/twAZLFU6eu7Nm3ln87RN4srPp7/XCxKMXBnV17MWr4Y/B
VUzPpFpnBHFOGvZ+xlKXneBqJb8ukDvO5LbELumSSbAvqINHm9g3hg1HH7Hh71hVsNtjlS6sV7Oj
zquIt6z2CCcnZBtg15yYmxeS+5OeMUZvE2E8PWZGdhwmObXPjhFk1W/CYxf5OO3tYhdBCLdPzh4w
/4K7oznyPTRERFIyOIIXdyycAiGO+LJNHyPxs3ECBEdqA1Ck67ISIA8+NMETtd6OhSnZ/ZdGbnAA
A+/3OS3jhuHHGfw33zmncJ5Fm7xTAb45RussIUPSD096oskD2Xog0sAZRNGIkMp/PWclptEUWwoU
nEl7d4n25ETXjv/qtZwp2T6cU4Pl4e7AbcJ0+Rk4aZ7A6LLR8FLFtfqgdRvhUN7gx5U5CdHZjfAO
BSAcx2tzo0piGAwtodFPEAi45BvXrsRD9AKzfhihMZLF0C6Pr9XKLO5FJkC0Jdr2e5awUHlwkcts
uZWqSbc6FlrKbsguUW0q7mMki4PNqptYwzzPgSV5ua+cFu41LXwm2XjVZPTkIkGsJoQCe0ju1nII
yC7mw6rs10wTTlMWo9JU31SEEycO3MAKP25EFCJlGEgDeuUoibRzsMtsSvGjmuZatXgIc5rjNmV6
zbfHC/4IPdvsg/eNVNFIzqWX3kySMzlUDXB5igJGK1uYfGOHfa5Mfr1fqwgCXK5gBDb7CArANtur
jbUpXjDd8r6KhJdegau4M/JkonTkMwAmaW2uN2lkz7YVS22XI/XlUHSJZWM6PsKvQBmbVwEEOnSG
cNnejQ83t8Vn0rRsV5WNpgmm2gr8j4c2bJDHUPflimQ7gD0Iecz1pRf14FYBkk2iH5sLb5k3ldFU
8e8cf5Us3jIPJJXDEvtS3rTF2nbGez1KPqzIqzJnqOnW7NTiVZFYMR4ju7J45oqnlV7O7HR62GNu
FhPuhZz0OPNWi17uIkvCz2S9OcyTu4ZWwYsHQLSyOLg/6lcoiLMaivEgqOm5opys7pZVyXLdKFlg
Fc3B+JLZArAr4VrPivB1K4WVWpGQg0HrfyQ38YR04dm5FTUu27wQuW+z82fEYriir+PZPgv2OCYs
b63z8l6uINY8MMan0cKp6dUl1df+DBs07lBwfwC9ygtP8yJ3m6YizXWzfwoeS6Ny76AyMhvHy/Lw
okoe8yVmQRBDM7SvwyUwBtcbGShrsjq64iTbMkM+xizB3cKAgVOrw3wIqBPFIfSefQg20a0AzcBK
asuZpKxHeS0GDPJDOgA/8f+d+CV/NaCUPOtey/NOI0Bq9UNaq2cUpfxMItW33BkZrSEsgVbFODN3
Q2RnsMsHbs47llasDrLomINuEb3yksk41uxYKc0cSvDicSficNl6fgk6KBSlKweFlDrerHOYK4V1
ADoiMgJoZ3SRTHGyxEIGZajxQylBOOz59UTn2O3bfHYZLDbViR4ZzRhz8EV59FOcH7QJcfF6ngcx
0H4BUMKUnfl4TPBUJGvbpKenL+lOekERGo/B/YSdFF4YDfW2oGgKtKaW3MjDH1qqRh8H/zW84R3/
vCdVrlDcCuPEhTFt4iGHIoub55q/uGfr9o/UbyqV1IL5uX8eRxukBVx1OVuVzHoLT0dWEAqFzLTN
ABa/gb8lzvNZU3RSqQvj9dI0nHavJ1bgPPKrlBoDixUXval/YDurFI6AQTvz6hR2fUlOOarExYg+
tYykup2dNmM9gO+AFuqtX/S5UFjjGI4M7SdWfvOQvZq6J/EaYpWTVpY/Bogc0yQ7mnSfXNeE405B
gP4lHw846akO1BPXzhNWD4PSMhHc3pm1Wl8dAhafIlx0AU9XrYBt1RcVBSEXhV8JEauV1XpXbxwG
sMtMLXB5CHS2RtyyJTg667XEtN+cdnvgUbE5ikmRYqtAp4rT8dXgu7jc5JavoVGRH2tCtSCdhd9X
ILTvq1hqJ8sWcmD5qLuxVwi45AvlowHS7N7wmEJ5cZiuDvbgN63cT2FWIfhKhkLjnFt5j6Bxd4Zh
LHCaYqVyA8djfefgoVasYXn556yNKHbpgmpjN5T/kr/SQgrslrth+3Vy/hpLHI1LIElh805Gl3oh
DyIZYqrUXURKpxOoscSKC9pHEroFbagHDzKnemWWNlU31e946RctfY4nxyHrLNCfC68r7aJOtmL9
OfQTD4w8pwBUKjTvnhINXuLw/wyOgUp6Xx4Ij7xTk/5gUipQKVSv0XSum9eRFmYMO6PFX2UtcfK4
9Mu/ZmbWu1GS+ckCRGJ15GWiypQbi7b7siOb+8QV9bRVgNXw8o95UZr5T0yIhnovANtDNBOc4Vsv
YFb6utqMadGfll+NQ0X4ECh2PJzHR/IRSwRZJoR5J4/eQNKIYr5cJe8sL9ZCotrb5SIlRJri24mY
pw++6KjvZB/juMNIWlcWKZ250V1MpCfDI/BrmOfsO5Lj8W7XZ4KEOQjG9sQPHWaqvATvYx/Y91bH
TsQgN5y+ftG9HBISuUXy7cuxqmcKGktvnet4jOwe2w1jsx+q84sDKk1dK3vyBbr87s4dENOfyaBT
MuBFm1sjNlT+C43ChOQ2fmJOR31xRzpbfbPR1EDjwYVzsaF+D0FMY4x/qpoogmsn56MLh8VD9DMt
txUdH2+o1m9BuWeeCG74hoB/4ZnleT+krsHq6HwbK9PxKRDWVhhTVhWeZf/454z+LtAHS0moEKSx
Sc4CEwO227wPgrCkDL1O7acq31UUEgZSwLIs+ELCeLmg1n9OEjgD4AnEoSv+UnF7M36++XS4RAxe
rqH93SLfspw8HMxlZfE5OBMd5yLbNvrdyp39begPGjWBNr2tX60bjhObaiqsq+tY2O7Ydbunt8h2
iUJdLy/KYk+mk0FRbQeNuhnZ2WIOAUoJNaiPG3PKb88dhBClH9NmrwxwQDqwtz4rHevBlr2uRI9C
4pItXGzvy1LoCXiGMEbRDOQ/3PkDN95jD3xfvOEAi0W/gikdutrY6Pu2kHw+WHpihPrPsStsQUN/
fO15gHWU7Dkg7mm3UvGlE8yfttm1lZ1sodS3oytogGySHd+Hl6dcBKGvNmMCvhsrEMapfIP0qvy/
eFV3XeTQ8/uBh7ayCnIHG24xqq0S43SnGL+bCiOjvFq+cc4FUjsKR4ijkEADUIYXturiB8XyMONU
vs4ox6i7c2bVCLvPaWn69h4FtCWnyPgFRikdTsOjrOK8x9Q/jD+Yfidg4u8FCXEQu7whcMlcZK3i
xJ0Wfw1YCHa3fDc7xN3K3vRNz+WkJ6DXTL0cfVJAPtF5re9ES1/ZyPcop5T6KihunclPu1T4Hizo
2Gx5DFliXyxOwySXRCch9uHEiwN9Bso+RIIcStk1amW8hu5wBetxwXZa+xTeixPZfMZISFqjYM1q
/nuNxxFocz87miHDWKltR1cNopcKvXDUOHt+u374R3TZaom+Iwfq6O4Ghz23RNBm5ce7orGw6AKr
EqFe541BecSoCNV3AGOeR8c/mUOXJgqnyH4IIavxcukHG7h6iXw2PDKAPkhWnYuFK/ObxCHOYrd/
56twGDjbC5Tn6UQTXqk32/kZ/iv9frRyP/FcLWEeUaubgFpO2E6e7Xx4m0fy0ND7BhozRA2VrdX5
8wQa9i4Um2sSQJ5nKyWt/9MzBZILuJdOXyfIyC5gowOqCJzvrp4Mm2RTNILUepfZFHu+oPOkcrDt
2TiL4m9rMk7p3tAjSOAy+Wp5O+go7pNHTaCRvfebuSVbt62fYnAagjkERqrkNQlmZyqZi/c26Wc+
cZjm2K5cIcXHZzhP7p4kc+14AXN+2wTvKkeQLiiR0Rt8aUjHcrazkyDZp1TcvM+Nu/Z8OeciA8j3
oIuCCKcTePEmiYaOe8nr9xtpkVnR29qnoTRmwDVs8xCZF7L9aH6ah02Ib049HcxA2fxjD0/L8b0Z
s1vQfdqs8R1k6/+ZFC8FT/IKJ6H1YURnhT5ujAFoBAH41uGM08j9iWFmgR4kQyxuV38SD7wxBQto
iLxzLftAQpBYbEf5ekSoHJ67gV7MUCc6ON7zgTm0W41kEQAQIHqGbqeMU3qxbAN+5ZewA1LxZDoW
6A2ZdWAab3Aqy3kc1E62hnfJhvNyP+HT8Qk51GtRoVPkZanbS5wxAo+lxj/VRJ2VderNXKP2MMc4
MATWK6rAOU+RPo08SoCrl2txS8PODlEkE3zbBFkUKyQISaPhEIZXI9eIVJV4BOG969X6ugzdPU1v
rOfuLJRtFI527fHDnuSQ5uagrA/6O3AMT1NVFnvcd+yq7uLi5ppQqAyZuEqhDWTQ8UbYeGAefoJO
mkrnga2llwnAQyhsFhATUoLIvL0kmiYHzI4EXwxk4lrfbTEQw0u3NfVVLcFCwNkt6WqDvrDJX4eA
AIqzW4Bu+LRc7Osko7XImNWSZNros6EJ5i5epvc42bqVIm1wz+W+9vrhRrlI4n+3OGvTr7JxAvQa
yvTfJh6P+OJ0+BMHWA2Y5T464jgDHLO6tgDnOVx37rYRTifJu4ieELrGSlqAsqNrMQN7di36QkGn
YA15N7EKASJo7VtCsAMRl+aa53HuqAP3O9zo7PYFc6Q8I9Af9ACZC1EmMsVoUctNIX730Hfk9ud7
iRDA9exo+fwLzN9ewbE7NXojSmQnV1QA/LZVcbMmwK4hrjJpL6N6RKmVMSaNbNkI7Xacw0z04CxV
oKZxCg92gdb8VnKoqfyIIxUG5DttMj9UcOb635ZjSVJS8XQArifIJc2xDTwBNc54pPWPuikKq4RL
QffBqbzMo5/LqV3oRHIc/tceMs4IrX2dES2cJ1WzcM4HKaDQNSKq0JsPSGlUOVMaWdQidw/Upu06
Y57v2F+HBvfi+4gNFq1Uj2csLsyvxnIDmI4D37bV7htAG7QT15uesos41TJAUfxlWFbUUSiwYUNC
G5Yrh6c+n90K03PLRARy/h08l8/CxYDyrIhvByAcExkfxzRtP/t59KU9F2F5bG/u6t4rzUH6JKrr
E0g7NiI8xi1dqwgzzzjbFcpnvSQ/yTpKbni5rXVUzXyD8L+vHieCGpPc2cxvC9WDCH1CthZ4bAls
rC6f5miyN7CVc3Ungrjk+UHJvYeqJF7pXMNCpTFURHVMXeTI7hVppRJWyw0JJrHtA4kNwObbdwvR
GfmH/4XbRZsXjI7NdL3oMC+wtjWXZ2NspolC4tpHrNk4uR33sC2og39WaOTv+BWW5kpYRPXzHx7+
G7Q5Fhi4A/so/8WmNfcqo9xPeGRSygB0rKUcU0dp9YRblKCa/u2tazvXw/j/8jRSwOAJT/GFvBbr
MKT1i76R57XBZRI9pRZ5aazOUf5vDPsVKXZtt+6XM1u5eDfv/RoATbIoKN53TVuei68XWAU+0ieU
DRVprKkxiEu4gNKIm/p47G9NxIfruPiizahqI8dARfY1d9RAkhLP+EhXz3IH6LGDxVhAx0fVdxg6
ibqnzkD6mByTQQBaAcxzIu26t4t4HwwIOO2OQ6o+y8YXaaC1i26PkzbbGnMnES679iWtEa//Xn8E
qmvLY7VUVz4g5VtZwuEdd5cj8XJPbywJyVG2xowFkwE3EgtgOfaHBk5Ghz9iTISxjRVHoYf8K2SV
I4ZiQ8aZLVYMbPv7f57dgJdYP+rgbx6ekKLn+SinarbLNNZ8WzpRcu08T2nRTfy6D7eWvFX8oggr
fQo4L7hpJtWy79ggbeG0GrtYKFMkP7AkQQmC3St9CBpeyh27klfZedvrM8vsKP3cHgqRLZQGF5b4
UoULFg6s/ekK//ZRWQ47mrcwuPH8wHZRrzrwG72nsau6pQH9/BU2i3NjMcjLiTCBP/dE3wumItN6
vgCdJ+F1r545p/dS68X/M0O9V0WKEjdJSd0J3LigVwgV0KyNTYP+K2/v5ViOtRNDx8Rt7UuQx2OP
kHCFr6M5FstpMv0SQXrlIL7TJuVQfCLWFpqJ+tvPWJVLk0dck5LU/LtM6n99HS6PvvJ9dVqkiSXU
6w509+JIr8iKD8YbekhNeDEW0vfA8fSBrLvLkSCRuyex2WUffgt9R1cTqITBR6YkgOdJ8dkEHk45
j7VN7fR5a6MWl+0AlVQyLn4cv70wEu3+3IAZl9hsEvhBEvzhKgfmw4fSooTXUaaqXlh2JAJ2EFZY
Nf76uoYVakSvB7Y+JbC61kNns9/X+g/Oc1iw7vMRSDUeIOK5MwoHIm7/hrF4I4cp8Iu+cRZPPBkR
Yv33XTF808hhJmm8LBb7X1uiOVWFtOFCTTCsOEcAK2QN3kB53jgSQ2B8hXdz2nOAzNeTAD20lkir
Ij4nB3n4nAan8MkLJ7TNP8fOlpeDbSjzqUup02f+ukp7RRARmfSATN++cwPeodiBPuOmkavvi6oT
QBw5+RaaaULBnjdS9YHmpdOuAZ81wwjLE9dkTXXD/fVpnuP0zxo6mqSlxBH2hQnIzfm6uxaHf28O
J+Vkmt4IZpmp6hHk8Yu9MZXMgqNkFRHyZ3gtF5dMsKGAOWdSjfHIbKP7O6hzzhy3OHPGwjZU8bdq
44H7MIEsqjviT+Nt7pfJqzkKQk3M0yzlBA9LCZzJAR+T+eZtjq+lmm1OSL51LTmKGOVc5lj/Jgzw
5t4yuz1hYlBcSZ/GOx1PesQQ+IQT2g3dIQ7956nzSG7RN8i2aVVbQg3JxT0KKAreYq5+GGKRrxnU
7Kv/qwQBnQNg/HYWx2MoX9Kidr6InsIS+4aRtQAQVSv61VGSDhp3xKDmNOWMClB++nXSdUCLJJ5w
NH3LES5Eb7N1msACki67kElzBQhyfaP5gGO3wiGPYY+hsF8wjyydRuXr0ImtEkYldhL1gPSdO6x1
Xg+jfJpLYdsaF7BaLeII7YyCkPnVB6h0b5A6tPUOPZCIvl6MdmJRmjuCpPwXzFqyd7vNGmuT+Uvg
C2neIYZDeOdehNk+dWWfgryZ5T2SAxOdz6lmVKjQVzcVrhGJATSyB2anhfEy+0al4xxbdT/wR7Q1
N37jfVFHpM/d9IL6lnfISdU6sSnJHlHMkeoHSFShmmNh+lICbVHniTwSoJz1DInHhlNcq81xp54R
oFqR/uLVbzFqIguHToYEjDqE9sa/YlKQCESC3xHDkY8ioP27RiudcEG2j63PRJ5KwuOuxPacuMwF
2R7/T5V2PD5KK+TujNprrplli+EjQncboLwPjurUVaQGkBttIIcI3VS2o8RdMtmAdatniUwJnhhV
VVv5llOr1vFDNUjW97mdZV2/h+xjgsf/UtHHksfhX0sJI/aQ0Ql1JAsA5u/DZf3vA7aoeNYfUtNE
sAO4MHM4vlGc6o5BJuKhjgXWk7I13KsyFLdGYQSVhLfb5v6/aRPaVKEZb1rldo0RuCAmgHnLrDB4
HmiBd4qY/QiGsFVmwBKvP9g6DuUrXlPMHf5EIHy5L/5YAQL33ABO7J8MEATHDV6Hx0F79RqvVUy5
q+3qzwHalWAHw/Bh0eUdgvu0cNEYTsuR4h0QdMMkTekZBj5wzebjGP0FCRRkwRVIa3577dVph2Q8
5shj/iIsTWuCI5Pq5sZoBoi2do6Xg2ojdF0qsbnReKjzcehqcH5kzZYr62Qzk/husXhCXEUCwd2Y
00CbvM22S0DC0Ay9CY18eISgRGLNL4m0pDdlj6KLkEW5YMdJhBDvi5D6PLDUqDo+J7ZbflkdlcKT
wYMbse7yFqTmKJZ9Y666QR0OK1D1LGok+nQXwn5bWR0q541Aa8jTJQPbPQR3A2KIBN4eIpImBmw1
MDfhmaBf6hvJmWMoRe+4GDLDhxeJUMwJWajliHSgflePcD4ctuTc1msRHxXdhW5Hk6AEvWQyKwWe
QZ615mUEOkHPISXkqKP3QEfong+R3uFDnDaMTwBRb+eR2u9NdjNua4kw1iHQullGU7lC2Nbbp5er
halyaTsZA29+YtXLqcvukaufX/DCb+zAZe6GxeP6zRlu9qzJk4+DDEcbUu7D36od3lATawakk4/r
iw3uy33dstnr17uu8IGmyAXiWa5YB1EiO/igEwny9qPpmhLUPfgp0VBZ6FIt/rTT71RMAXr0fwA6
bG84fL1iw+a3zQbit/vydT+qOsG0iRt8gDzjeAbcXF0os3cPrFgJFX11UlFjCiZeQctKxUOWKBKQ
Ulb8Uh4RXmyR3ODCx8uQBzhxaK3uc5AtbOzLFalWub1El5XDJNwAW0+9CWu8dgZNYybCG955D5W3
Al6YYf7JSpqaQkyk+gCxuUD3/gxdml2imDQPK/kXsfPU2tHBUcrU77g3pKP0UkJcf9xgk5hpR2M2
mCgVqquC+jZE8afTFFuR9WmMqjgp25yW9RfB6jhrnqvxHWQ2PSD6rTBf0IobzYCXnnw6wndxzqfp
hEGuXpSGUpdFxBBgS4zd5wS5Z7+5FCn5u6YpPAMvyla3ckXLHjJzFMH25cmvbh8cWlaUoV/AFkb5
DDB26j43NQjmP5Qu+yiqQh3FCPh05elf/hJmlCiG1YcMVqu558Sz37sL7UiD57/lUPZjJO0LELEZ
r+IBg9f9kowuKHNeYcE7bj4HOXlsVfBm1Kj7mwle8s6Pt7vrN0BvX2NubmNcUwjnisDltdSZDEuL
KLot+UJMzAlPSl3NZ48BsdhYPglexlX8g7pDkZcOwQcs9hW6TYTZ3LXhMS6FvzBKfm8HbvRLJOCa
NW8fkbQvDgE+VcKSIJrC8gRWTu4c7uuKkM8MEKdll0x7A+Gnd60pbjGi6igwiyHcIjycsFbDPOFe
kKVvf33o/rAUCt8F0nDE8R2KQ2QF0abSqVueuFP2MWm7DkAftP2LL1ZgR6g4MdtvLuNAItLQaJeH
MFiqd9fjLwySMk/wQwzqAxLRHHvs106eqwqGykrxTlGqi0xgtJGFDtp0EUzhmoAc7cNA4iFFf8O9
7x/F4O8tVDFzMelAKT6teY/ELXy78akTI0j07pAunxWpjfrk3i3VKwbPkGUC7xd6kx/qLOEGdTkk
lR+01sTvH00tILl27jwFuVeVXRKxRgAAA8UdpKWeYgqrfFnbbrP0NpjPn81VSxV5SsemE7fwq+V3
rbGVl7sbhiFipFThJbDILqmzhClh4VpaZVFysRmIfBa+9Od7Ja/dLRpZ3Ih3k+Fuw53OtqQFurTj
reVEbsfwbFXFopAG9rVPLtZSoLereCcDhllT6srwVi9y5KZddNnVAPCbmadbcw/BmL7pnRNPqj1k
e2A2VsbM8Ss1NUFnSZW+CZHUI/rOkm9YEkLs5PUetrtUCwwww4DsWQ8rgwzi72KFzf5jULl1JulJ
BblwMaUUcs7vAv7nOD4S6KYj2/NRo07gsCO81HpPrKAEJAsH/OkDb1Bij91rbqBGbvLvvchB5UjV
Zi/nBNFWic3cF8ZHkKH0w9DyAlHQhvuLxc9pXtc5OXFxT2YcIxHHostxBKHnkS6t3aAtmyJzaL1Y
PlGXB2wpDoQFoiXaFJodAkVbzS3Wcob9UcWsuyaXK8VBnnNDLsUFLMZyfucwCWoYe1/kBbUV1bUW
ihUXwKJ9XToG9/3S0gpsHtpd682qXG7853G2jSMcvvd4lVMlD5x6fqOx5J4/IQP7C2njdAKGZd3D
ZnaShKSsSOTApSJxbMV5+H1q0TroojrRbwjMXsU0E3KuhktY1N9h1YCbZ9iBh1Q5eT+nAvkitS0V
KeEfdxgRipfkfIlOy4mN8IVHu0M6saGGockUKq3504adjEA4m+FjDbSFicGkJnEH+NNQU7oG0TxJ
jUIgpep1HdEYkvXt5haNn8kHYPFcYE/8myxAxRGEI9D/0nlEYoJ6TbzIy99Eiwj3XkTyqFy9pKXp
+3ycoEwtLrQoCIVSpVcKEVWvbhb8VrOI/N8LqiEA13APyhfZh46NNNutT4/MIusEJ8NdpCEI9VTD
yjme300VSltGU411oclzRG/DKbkjQWP7xoxaY+HZlEdS/vjNuKuWL2QfSANJbDOglv3ykNRhoifj
14DiJNkfGeYUqzGbsjC2s+p+HMw9fY8TKrch5R4+S7tctyKw0zuq9/oAlBRuer37A1y287iNUtsn
nP3ZBYsfYzvbPDTBcblQU4aS59BfTtiSHsYmbvgUngcqyKCfiKJ0PD9Nr9bbYhBEPYEbm8YZMQeO
CCY2Xx3xLNTTOQ4X05XLknrsEWC6Dht0v8gmq1eCtoK51GggJj0ltzJLD1kqYnnHWaHJPGOzOtXX
6Cf+9COIYAYLpuHBoMqVJW1t1cn7WBxQyEowbBTlfeFXeZ6ogRXtkn3lVhPIhWxnUxTlqH5avQVZ
bnm0qml+5jKH+9JJtDgOEFjuUExZuWMtYAMRigk5wGhrYhTjnLm2JNb0IfiGuQmkebmnVv0oCiP2
FS1rs4t1mDwEReKGV+imLz3hS3BizyW1NDX0oUEknp6lbRygk0gioZ2Z/a+1zmDdCJf37k8cSq/b
5VgdTwkQHFbxgpzOKkhgvArnaFK55/+TLHCUMB1corcfeM3qi5MKVEl6j/Kuos3jmpNLvoRDz/g8
KaLqQ+rIx1ZDrTf6hXvsf1iHjZQpWf03NXvPgSLxOuPEg7DuX4GOpwBVdELCjL1S8ZVBRw7B3Yq4
aWaGAfoFipjaRvk0bmoG8urUTCBog0UsR+JKeZFEvL4NJvB9tFxYUMmQgbBA1Zt/ufhxFzkDab4c
+5pLk2Z2x+hc5S/gu4lS1KZ4c8FBhmFxYGjrWJDAJygrz+TDC8AzIhilT0gBJfi1fdZeGWywONwH
GYAmMC7Bs8SY42eFnoiSQfWwnQ9dKSUe7UOj5c2ikOeFnXKReYDO/7UyWlA5ONXxQGBQ/zhGu5V5
Z6HBP7SUb1xweMj1Sk+G+Rk2aVehkyJ9FfXBlYF6C89/q8gmz0XDu+95dMqJFjU+Pf56nsyf1BtM
ZVidK+LyhDwj0oYwN7C4E9zKacUtZZsFdzX35JIlYnCGfCiTAAMrhVKVcZH6+6dkL6DhuZlJ6Cnc
lWva1BIdE70h4JCILhiCuEePBofqTtZB6zOV/3D8u20iPowdzna0smlqxqk/7vFKgbX33f2P7i31
1BfQKaHRizELGFAEtws7I4251ovCr76+pTshJRLE0xMqgj1pgrJjRa0DYDjWtWMHIqkiddzvxhGc
CrTl0ksv2ef+D4gyJXmYWgfLQBJofvItxUBEXPH53U2ZJN9atGEYC80BoPcsVXF7v7/b85tYUHWl
Opw+R26+0cOt2mp47nDfziopTRlQYMWYzHMFvauVjaaVBcwQnC/xfpXMTl/l59eAeBdkWwv9mRwO
DTiCBEI6VnJdXhX3h2YVV7+qmZintooO5nGAq03KViEBK01mit5nUz8dl/4pZ6Y/V3sbPL4adgCG
0EUaaW6BGaxk7tamiVboyUZVivEL1+isa2GJJNOE29tCA9JZwTkRDtw2j46Jb1rmZ7q82SDPRFBg
Ks35A+kbobKxrKvy1N/XcDXpj1KtEfKr9b1gFTorM5vpDxH5iSIQ/stG+XW85WQcDWNH3MM7bPxT
sjBlJwGTyLJZxne9q+4VJD0Ew87ZKsl29IRRzN/PMw/pXYPp5im4HfnuJWRhlI3/jrLFmhm/jDSC
Rmxx6DXHW141ecEregXPZYum89ewpp9PJVB+iTv2A0HVxNgAdLNs0GEf1ynFVdO/KdiACPSQMvAw
aT7wHQb5barv+zHLvzINmbDe7iezdukkXGsb1VHa8mXtr3pqf4D4hB4VrK8RBYNdbpwhkKhNtp4c
p1MK74TsTqHf5gZxO43R7TRcy2t+wBzso3MZmpJTRkEkSKmPYpy2MPXTgJ3MfhgvLgyZ+sBXKDo1
7Ewr0K1cYxuXwBQq/8+qfn/2nXtPPn8/1qDrXvj5doAFcGgGDaepE0eqX6f4xQ9Q/8EcNImERaUE
vnmFkSGD5R2JNYWw5Qif6K8oOktd9mIioViW+QzD+icaVkJ28nmvjO2nSOJuHjEbtg45+0NPCZJa
IUvORLUbRPjK5Smv4BS5iQZ3okIJtxQV8kRPSrPcO+d8GjMDVIeaIw4IKaPyJj5LcoNNR3HDZx1j
nnaRQRqYuPvi6bVkb3c5S0EV8m+Q1mZQWKjA/WbHOsI56D/Be9uhk0zyjCmlErAOMjN0P6glJPYc
Q4yytadCDDGR6DGUoMF+t7a+4Pg0BAwN4K/yrhzJfg0EnSTPdxbOdZUYJ04J40UrDkrgHRLeCRxD
K0KPWv37Krxo6i99stAa3H9hwyBOxn4fS93OYN5a3Emynat/6xApuxhrcat0QvCWg0YpNAB9I/yg
NVfRHmKrlju/uMRpS+l280e17mYHZZW3JQ9jWm/CyMzDV8qbeoVpI/S/G5xTUajuK2RTRyBi5R21
8krXbVkidMr++VylLR1jmQ+YSPgF0YxalZ5i9ubt4M0r7wlsp1xxMR7O2tiVpAqniAcwnu1veoPA
YVI3aE9W8XmntD31PrmXOgtF2Mz93+VUYZK83aXwEsnpSSyJvdPMFaBiKZdhNy+6qhRVFs3uo+a1
4HkfKKTYT2G5smWllYBblvVpdWF+r5dFp5mvIX9LztynU0CEN5t67q6L7xkcLC6ruI4zKRUvLbVa
B8kIUL5NBfdeh36DSDE+5znudpZcCMwVJpMtLVSz+VEDEqgsAVpB3UdW5RsOzwJ/LgNVsS1REIh9
QjmhJ0QL7sYP/OXHh+nODU1uQlIY2Ve0QBiahwjcDzLrqcgzn+V6cd5la1EF1PPYJAEOZoKJTina
mXKJqr4jS7PLqwgrMmeNuc5bSqsbfciH2AStcTifxSCqLAXLlrpTdgcQzUeFsL5uagbM4kFMHQ8G
HqoP3FSFx8QpP6IoNdDGMtz5jCXAIeCGOi23xQ71ecX42QiSdi0Io5hmJy/gG0fYrKJfyjUQEvZL
MjNnop1fNHTsB4X4A+rqwIyaErLnfJK8mFYA5saL6UBhefioj2Q64Hg9bpSj5ZoowG2syUBIxXn6
5wd7YrnED/RmUhnb+iarSIvHszFaX2WC6v8OUAn/MHxtGccDw58JTpUdjJs05lKllX9DBCL8yd7c
bd1Acx6v96FqCzWjSx7KB566n20dUwIPhButYcKhUpXSY4ERexPCzWNH60w49+de5BDwZowQkvQ9
Z3X8sxYiJ07k7fRXFkj78O7X8kPCbW+Dci8XZqiBqdeqKDb9iso+X8kBB0SS/LNryGTULtXm/FMr
kN29eoi4ZquqYCCPT/9Cg69+1fECadxdzxKdu3AFcSscPLjR6jbzxhaEV4dFV6yEU5z4gRP1M6Z8
pBaHsyvor8G5O0FyDzWDf9wtqVtNRRdSoPIJzhSHHS2BGtK22g663K8Z2mJSVZOfJIW4SzWU76sC
zyhprmSNY5V2WHklG3K9/on6aYAmVYCSmY9dGrjZcSQGsUACb191M/pjpI2I4HOlxtaEdfaG9K/E
/zSEBt9vRkGGQbcq22jpegyViIq+UNKuZxaKZVj4JslKc+it0BsEhTM5fQjHxy04RBtA4BMiyRua
J6szD8GRhX4LAWNlJCctPghVtEXac9mdq1oxJkSeqspLspgbD0jTwHrnxX7FBf2AMOCv2apLXHV0
EK/Ql9hNGGCsUC+G3CzBuDukAEiBeM8XnrJQDGqJ4Q5vc/C+IR2PMsYPj06CjZ47NCLSL1DnqIdM
m4hB8OcTCz27FhfQI52k/pmYzLnGPBiu4wP8GstWZpoX9tNqnBb/RGbKU2+w8hbbq5cOcFZiel2r
vdEXQxLFQ4N7uNNxG/od/cv1VnQtEgugCYR+flJVuoqYTccQu9HMTUuehY1hw8FvEnYW0utoItn8
+Uf0J74Cn13AxuiaiVyUYPGgQaWtAntygbSZwP8wOg/2yPr7/nBdyXz1i5B5gmyiGCVyAfbbrA4y
WMptMpfRgLDIh0FW85ed/DDplslN/uTg9XzDaCET4OKqUbKnG2hfN9otkO3okaKocZnz+oQ1QNgP
Y8HXivCSTVl4U+RkAPI8HeyjqWjc8swx51S8j95wQUw/q7hTkezSvtJ4lWm+pfB+03ROQDQWTBlI
C89LryZaUvHsIm+YUjyV6jqhU8JZRkVDeEr2OCZfF7/loK2JLju2jtMoCrSyiCegqfe23DBREvlW
4X1wt7R5yPyKb+HXlprjhCF7BaWer8ee+VMPEk9ZKugh6Gft3JlkB6o+Oz9hMgdLUFImrsHcltUP
oR7Ke6uLQtyQ33sO2a6Q7ODliNDOp3/Nv7WH7IuSI7iMdFvdHHAGeIdXhaSsdxvnlCQ/RMNAEiwz
dW2EocjGxZfoQE+whMw4DMlPaQKmbvs4/4C59DiKlVxSwr4d7QY5v4OU/GuU3c1P9a6tOKa93VGU
HsPv1HlspjjCEdSnbQ/0mbaisf10EhvuclOhh16dG7KtINBJGLhE/eywuMQTV/zobDk+s1mInBvK
xnTCGWe2L547yjKWGtdrsNGAs+cRwnzGApBtyDaezb83wIZDOV9DXXOBIYlrd1MqnAgn8TX+Oepz
8W3KeQdEDjJ+Z23bpPxgv4C75p6D79Cq43dI3cFHVRLxS8ZOM0PQ/YCXaS6U03wEb3AdJyTzljQl
oSGUz7FLI4MRIdnIWRp0tFZp8GJ3V33EmIOrTqvsrzx/uhBwwa2yHBVPP/eYuIHVYYFMLPi/5+nw
t4pRJoY5DilhGkKnNzFH8MZ1EwO0zK6ab44KKExpDo8LZcbmxvQfC8r3NXMUiMiCmakCNtZ4gDsZ
Kg+inRGNSz1dgcTNWdzoGWFN1IG5oA+0DWp0B000aClkrbmhZ81+Yt+ZvZgh4wrEGdpoMXmhLCzG
nxCsLs/85OKoEInDZXL5oR2L9idhF5wAXBfDmmurfxw/525QEXG8pwGk5VllZnbw48z9z9mZa5io
JDbOoA6BE0rbcEm6aUZnh4WQ1aKz8H6H49+cW4YKljC+OhD9xIvaudbAbWJ72hHl0En4h6+dQMqD
F696GU1R+Nr15WwmvdpxhKCE8EM3j4x7Zzs/WWH5rVJqa8Lwt9/e9zOvI9hpsPO0OkMRqfgmPpj4
hLue2YYtL3zUDXMP+QGG8QGO9kfRU8aofihb3NgnNDNNa4RhCe03e/QfylWDPa59l55j5HBOjcHq
mC72x4Hlq2FBPc0qDlXjA6XcOqrnPcKU25OfqUznEY6zb6tavDXItiJjgbFGkX9960MCZIqJZWUd
wEN8GLTVclfJx+2lm/ucnPpcQ87sh7s+YWumMLd/F+kRLJxkeymPDYD9SpRBjxPr0OpHZMvb1FBa
nIPVreYbbR2aHC5OCxGR0urVUHP4EJKlPrbUwHEornAPz2RtYLjuGNnWBK/tXz2ahREl6MZfqutj
mASAvzIz4MpUnFzR24Em31t14UErktT/lZw/Jrs5ng2O4l1XEe0rJGorPpdTzg98or3+tX0KyeyG
UNW7/U1TP16QJhjSgmfLmR97hfrBj5+Cv9YOmLcNHH0Jr18dzXULdiGgdezc54C/xEGB+8KDpHLA
XZbu9/J7r1CxcntV6FIBscUq82hs3tPiBZRJTjzwwIaS+SA0TgDRVX9br6Ye4PLUxS6TpVtYD6iH
dwMhwjKhNSTrgHj5c5LuCUpT7RiKAhHtesdlNO/skOs97LrFBkFR/JhbBYctQjOQ/Q8Ta3f2Cqo2
pJ5ohI3BdJuu8c9jFwKHiOgGOOccMs4L5rsXEqtFEg7beGnNPi2AIBhTbynsUN6cT3ETPAo9w+Lx
vU72gnMMiFXgt4gb06srGZEuNrOMWInVSw18io0COxvSrc3WPTUh9NeLMebjNpc8PaqbQiDJ22oI
SWAHj6cZEfuQV8RRYV12B9niQEUWnc6cEGD+UsuMPI0p4WxyAsacKHqcbRQT1PMyKXSR31WBq3Gg
GyI/91qGb6/qztJW+bkrQvdtbNljyVG/d0B+LE3NoJgKtp2FF79NpXq7jDA3gJ0jxeSPOsxGyqz/
sgZeRs7ZHKGeZtEr9JcVLPQuqu1mSTl32o61ZtALJR0Sb5lIhrWY7lCmzz/sisS2VsXHrkZjewJI
bgsobRB9DFD1QimYE33G3Tnt14F4Tzc5tynVe6SU5lLAARQZDoUofdFmLwuGThoM8/TGb3lihIkN
c8Eby52vLhnXd7bWbD7S0MtDglTEhg6iVS26fCHUQjMJKLOOkavkcn7gF7rP79SQU+0kYvCyt1QX
qIsjb8SxFXZu1rVCeR8MtBtjV1mxnSlkBY6s5Mq+vhdlM6AQM0EgfPCc2YCfTKnWs4qgzQgNlH51
Ro5VO8eqPdmrp5YhHTF2fSPwUVv01duiZdhFKTwAfhaQ4aK05qUHgcrDcAI4KeFiNOy/M8NQm/mW
6kf4/qe5jGNEweMzpfzhZeLbK6gHetMVE35mqxxD7YpCSb8t3lfvshcv5OSQhh8L+zvBFLu5/TL6
qo+YTZgH5qVaNzJgyx8w48ZYF4cOw+FlpHyi67XbAPU+EHMMorPWnx3D2dlSQbXy60mfCFN0bH8n
rOnObtfjU+6dy4Zue5iSUJZU1Lu+RJRjrcOHaSUmM46ZeROuhH468YxjeX1Z5LPpwNkRktZ+x581
dvHKCT7E1mdTRGm8bBUK0kmPHeU0ZRMvUh0ekqDs/YRzJLQNV5hqT91gBidOovSefmstn89jNVOe
q7yBgkIslRi7A4LijsS34v+EiSY3YBM9MD/XJ17OPtL2QrLo1sI5QdAUJtWRDwY99jQ4DNu3Wd66
gBQypOW8ONXnddI36aqMMrWpBg4g6cH/gG/jBwIJgWnwlhRbt46LaaU09opoj+BdtZUq9AuRv0zc
xVuJjOgXDsaa80bEPoQyAjlNtm+fiqgr+74Sdf/Am5pUJdHgcuSng89i7rOUcyhq9c/5+ToVBVQw
eVVK62bE1RyKprsl00s5H1wyq6yt1dG04LWErBbneXwgyEihvKzzB9NK58Kp9sZMVLQpIy5DqDyM
xu6ecQ8uFdKeXICHuHYeqBEFT/CKvnjrUv8SEwTEepB4/brLFkkRRSE8nUdZFGwZOxdOkGlzwOUV
pjKdHZuNLXqUiUBLRCmu4A+1CECtaPRpLyCUj1IcVn3DjxqWb4zqLr4hHM602cv/ENYBMAWzXbu0
vj3GYHnomYW/xZLWdQ3VuIPpuF4WTBTg5YgsKwlgYdnLAn13DRAmR0FX8vO1ykI5G90Cb7moFoI3
UF1g4R06GuwX5w+GclBs9crTbiR40HaFMfuUmKO047WPuqq1lx7uWqJtl63t6tR9GqEVrxRd/nig
qbGxn3jsGMWxmtEeAbtRoouseuZsgAyiAq7TosCvipkUB33tgmUAF0e4GQ9Cll6+nwwn7MUxboey
NyiAHbpoxfOmBm3VAlQWlUz8Hq81FuWTyebd9HJxvDBeOuJ4Dy3+6S0J8581pIxzyhefw2n9Lzie
T8IBZ2HpJdwuuRaJFALhRiwuurOuOedYbIrSgWP9QkQqnzK52Jrf2Kinsjh/QWqRntYT2xeOw6S9
YwsuoSPD44MSjAuQrpYl+lXuRVj1EVhUxiIT1E+2/Xg+nIBOx5x8utv2rs60u9vKhW0CfYyxs3NJ
T4OOEnv/xeGoIsMT/FxKMbkey//ymm5sRLnOpJhbDeQetpj350bAxwt2GZuZePQxjtvEliOs12/Y
N9fR9qF0IzHpxms4ng+yPdJEWONzMRg4vTWr5NI9S1Th9nEgAbt5g0WczjpTA6Bn1F3Dy5XKyQSc
3wf1v+1BcRSuhYWZ3nwla7d4aQ/fcCzYwpJG8ARVvCkRswmGKOWeQCeWiPHiHi21Dpgl86egqb3B
rzRFe/Ww5kaTn8SkfDH7DIXUTyRizVfyG3oct9DWxFM7nWcqWmQuw9TfJAPXfNnGGIZYQoh5Wev7
X5S1+M4dNGJs5yYCqc0Y5if+sh6tiWB0By90RvGpsuY2yvHFMciot+glCpvCnyeYougmHT9NRh89
fXPfDDCzbz3jttiiSBXwsIX0CYfkxPs9bPldTcY/BnmVNEpgcIb0M/XwwaKDjwbmQQyhQv4MI6FQ
vwMAtl0zGzxSANObmlClUe2Gt6h1Slrh4yNGInUU8pnkBZcsa2xT+77IILfxjswocb3tUHjxCuG3
Q+Flk8QZzm9uf5+Kleoa12xS/9FTXyQ0OKIo7OzMGJf+D2pkwbzgvo6fjQHnEd8rk3cuhckCoM8W
vIgVAkxUZG6j8XVIGo1LhHPwFvYI200Lqx+FzJc5LZ5x1wL23uJj26ukpods87ZcBw3nu4WYRvS+
ZulP9QP1VGXFMdEtjdaO9NnUwDtZARzLGMgZMidOoJbi3hszL0MVJT3Z4729wmo5VO612B1RDvIm
sHr34H7Q7Cctjig4/Caa0IpThxykiqy0TymGVK3zspiKpqcQjX5BFuL2Oi7ifzhRCScIaONj2D1B
f/oAF35u7bjtSnJu17Addps4NW81UlL8tz87ekKIyDBEeAbIeQnQSSZ6+IvxglmnMpuOga4LJaIJ
HfyY1TCh0OJkT1bAKNmqEelm5m7w0hp+bWp7PsnnWHGghH2epH+TzJoGkGk/YH54yirIacPnLZp3
DZ7FkfijwAg7ao/X/cFATUHwFus55ZY6rmFQ5iW8flUSCSxFVonulzKXczWdWmkApel/43r9c7pE
Ogo+8CTXVnbfcnZd5X2DNJwVoDNmRtn3oheSLMXy2YIlwWkr2nnlZJLVq34hO8vd+/fWO6nps2bG
24YiQvkJTru84TH13HckZOoCV2tLI0L42BdNSJlRVlw6ILlpFJovJpnTZx2bOalU6DuKExV0mwU9
BwWuFgciH9LstIUhtqjIK96C/kMTA3ZSR/PpXp7VprzB7g8impHJ96JRFhsCs7FhTPwLOHIyq3vx
5DzWQrUF+3ObCqK6c85RYVJMjRx8+gedmh4kY231S9Lm6QyN1rTs1G1JAp0NBegaNS+vLAKEIXra
J0h7o7ry0D5f3r0AhM2B85eDvZqT/RtBaTvgfhJAcE5a24Wsm4ljscXfD/6PeFSRQIMQ0UvzweyV
lKoz2bVNH5/K0TGnJ7MjqHLg0kmIb93KTTOze737/6RYqBZQxl7t1XsOKhwew6GcKsIy2VI/ShCm
8FJmcr0dg7qarXBHLtrVgW0DwyjKiKi34OdQKGCunlbFmWhXAsrqEEQR46e1H2usQkupGu6/bVoV
kjky1kmhdz4r1jCnd5RzRHQSwIjk0JtoXpbWISzMcJwxWcZPXTBgl07IXt3HRFbS4gkSv5FwPuPc
sWv8GdqNv3A44sf+pUxvM2zNj9pa0fEaxb3/UJ8FLVC0P+8bEE51wKl58l/tXL/UG3CHAweOqNdG
Z2fUvCNzNQYr90tHh1SGjHfWuQhP751+ALcvXmcgjh4FbAXWb2UowJhQlKX6IyQGIgZCwxAaadyK
+tFv5E4+94Nl1VriAUg5LZMAJqotwxtVfH79J3rXIsKn/W8g0eURraqv+Srxl6+jgxvhJscQ8sYv
rZZ405mQvN2IYzf/1f+/dFGfld0TunB1xiiHmKSWy1WaJ5sWHWp6fdQTIeoLWVjDSZBj4tPxj+y0
faEBzLEo+nHFUVSV2yV0ThOop02TfWr6DCEvhj4sQ3apTYybcbhpT1x+sUNvtIXKgFAMd01F8Q0+
056jgpfSGDWd4ZGla6GfO2WGoQmP4UNbaAo5t2JuZ4QENZ+RXH5WOPQD03u7l6vEoiLUTOdBPvBm
+s3Lanhy9rPftKmrZCnvhaANRe+atnVMnmjoOVrTYerBWBy0frS3elgzyuHXvgpKlmbp6boXm+JK
rJRDdGwMf9CZEDa+WOQNHJO6ieIMzvLuuBtkhwl1wKbtqJRsjBKfetO1obSuiMI4cKzlZBXUhPYE
rZJByn1Z+tDnYrQVwRfZbX7iwnm1a0WtlTwor5SGyf5cID6zUEWAAiW7+JN2mdNfEcCRjdDuPKWA
sEUc1eNguT7XkhKfsfCyICoxW3TxDsLpHNJiqviaT5P85RWIdmperc9UlKiPMIJKU2VzDYM0GoNi
xYBcHXttnIWUUESOoh60QgcFfztQbyT3CXV0tHiiE+tCer7yubuuRjDqrU98l9HLP4iNP4Yagjbk
zWC/Y6pmAtmCvHLoPR+yv8JvWtW6757KQ3l9nW1b+RmYbusSKSylNoWmxnmudGOwY5PLkTcWrqWd
fgIAyyePLFYit1n8GXb6m+FuBnyANAMa8JUdvZRwA5mASjylGu+9HdfUZ2Fl3gqwqnzFBIRgsP5w
/rCqFu/jpW+t433HEmzAsUG0yGIWFBl1kkoi8vqiHEgtD74Gt6q7P6xD56ah4jj4QsUVL3bXRHgJ
1ClJEWm0QnfwaGRnFRRcgxuFG6Ml34Hv4n7QBxAzhFp8wuZ83P39HFPExeeXuBK/a1mtScKgXQat
YK5OgaYC/cGDCqE7p91jT9OmD0bfBhQcblTUeQy4XCpOiQ9yjosJOI6Mpfzh3GovSlJPgJRx5mWF
rrUm6o14w2HTH/od0UlZwtn/8MQ1xk2wMtmVOn6G8nZ58DIno7rs/n9pjATpY6mECtWMFckhgXhC
nBaHR1ahUQHBrDaSkaheFNOgEVGPMu0j0LBlUaRHHAynhPHt3UZf6uaSakR9hdtMt/YftLsbA4zb
xs29V73vhe5jyJL89jQPs4n7BYX9L42Uxr8rxUFfwEsezcSoZqBV1XpxR+Q+I9fUJ8eePY9vFJFc
XojFr3wbSft5O1COwUX/E06a9NXGAYSGZkd+izjfD5dmHykbZIJkoYcUqpKfo7Th4FbNaUOzuWA9
IEw/Bp0XvV/+0Cu3QvL3xSMESBqY6zV5L6AQbEOmsCp5FkXMCTv4uveEYQJGOguGnJ18RJKPOPWd
aACIVjjm/tW5CQSNYsiuh6aNW0FTtP4D84hHSOpdsen/padOXiEKNKs33bLgkgyBCJveJFiylBfp
i1ddm2xK3rHo6izfnlNr+fyYKus3DgmcvikOaM9wpaOCqnfUJuGi7lNt/R1gm9fBuWzeRzG2aYDY
Wfg5XtnjqaZ/2HV7nvGV3/tUSIXSqzKcbpKOWbYZ1UwzKVbcmBuKmIX4O7gxG6DpEQf0xklFfa+4
aKNsgATvJfFl9q9erJxR5yAP1qSR2yTqINkG8MTQLUzOgo1+f5zDRN66UKou48XxsrGa8AL5UVB+
rTlOujd4WFBKwNnQOPmK1OP8GgE8jTTpWTerlK4fE9DGdkoLIdNnL2sUJg17SK9cTJi8qAUpvFbX
nhs+GKbXkMTuSRsemmhjj6PWqwbmOO29U8SCUryaHr7N/evn2qZyFehDI1o/OgRXlOPK0/x63R2n
3BNMt0BsahdxRcY5Ks2GLKNoG3wREeenkgWyWGNbsidFfWYlJVyg28ORqlHyCoWNqPRYNryvQqdA
SXVN70mfDeM8vcnVQEx8DwWgPR0oWN3VjZi0C4Id/PW7PzNF6Z9hG4tMo038KPGRGYUAR1EKFLfE
e0wmpz7IH2I1ciJ+FD+tsT8n6i9EmAH7FwRySoRwXah29oam5aC2vjDQ2TfrI1hu2Ix5w5uBCgEa
PQD80LPdJ3o0gVaHkfox4urz3uNJZ07WU2vifPNKt823Ax5Cqbp60nNdfNqctPiZ/JVD1op3m0HA
iM135isd4V1rpVlvu3VG68LSgOCtX350PUADBgcbUKtGoeyFbEOir9OJ6jWu/yNmow6OfqDwlCdi
Pnu65Cnhl7tMwz58SU3fxQcwQsTq66kECipMSiVgsEf5ka+J/IL1LlCtXeybHrTpzObyFfkaa34k
K3Fr0ehAWL2KYdIZzobJsGCg52kf1d4rtAr1p1Ay9ZM3GvI1iCWR+nmBN63DrzejiMd+xgm8DuXP
S7bJLx3uEK6FcUSg+YRH54apDR40iHWcSNdsxd2/c1yyp2DHoC5qLgHRJEeFFL8RIn5VLPZDRYvL
1q0u+1AimJW7bydVRUNnW5q4w9ClA2CShIF9FomTJ1EKOrtINDYOObKl/THAffFmorYAV/iYVuTo
mgJk8STQwDSsxfKZQerTcIZQpOD357iT1QLal7M/bNtzXskb2MwefXd6mMJnsc5x2nAPLCy7ThY0
GYFcul9FJDPiADirJKadvzytwUDsD+XpE1QMUdkPVvgsNVeWbRvUeidTNY9kC++i/dzej1yxTnYK
8iJcnWJSt1BytJr7TMDBLuAlSrki8gKiPysf6A6xduljRzRCtNOqk9h64QHYheAcYoP8h0kopfQC
bwrmK5PMvETiBMYyutGTBK4yRRWNehqzf6y2p3eGBmxPmrjObRjCQ7xJf9DP5f38+houb4pRgciR
rGEDBSmjnPeD/FALgqYCeXkU2Ce1uJbGGkSslQJj9DlmK5kt/mGAAPiqrSigtJiqvqyRvsRbUjTR
zNDgTGodUepmY8JcgWDyTbIxcdNxn3r/Y4NzA6FIsdEAmIKKgZV8ekgwWYfLugcM0fPXkuQ2nmik
hCDqL5yvjQvsY2DyNLITMHdeQL44Nait1V32C0fP6peSz9+yCBFjXZRUagKECgBfv9rmRRlYFk12
yqTtkGlVmdFu78kX8IT3mwhEQVeijbNTNoMfKneem6MuzGNRIiMruAaBra/vUACsYcTNYqfw531J
IIgspgvYiH+ce0LOU2CThgeapt/qRFPDwR5KsD6WNXG/+14EmhPd2OnLlMKTkYafzp8SHaGpoUEz
/QNpWQ0m3/cF6NMnvLOD27hVwqIzIynunk2b6eecSQ7WdsrTooDCS4pqDNcMie/ufyVgXIgKTcCK
LAeMvvjyorlFg4r9+gHhikhwr6WfxinKvENuOn5o4h/ef4zqrztxlmytgUNK6W3RcpAd1HmzZere
9HvP4khAn+wnhWY1ZQPFKLOUPhjeP1iuF55JZRUHVoDWrr2JgtXWzNfIGUdtCbHK1p4sXLWTthhI
tcc6xjgIwLreXuNyhlSfJI/QNa3cky6JtT6UTBuu1XsGfJLTvvPoZeI50TvHEhdTILdDyBCRaUGY
EUrfbBdJ8F2Xb6BbBLoxt8HtjSr2Sa36CZk8Qsj6Yma6ajU0DTbpE8CXqkXbcCNAQZOD0VDSLBgY
sXyl7oOicDIyHvAaJHcoqbOyq/Mp2NTwewowuq0Iezrivpu2KlrNBkEU3vFwYiHOhqOvhVMjGQet
fd04/2q1+4zuCbNLhMlvJcInODUHOn8/hgfHHvbMl1nyQwjMiXzNDUnFaEPtJZaZnQvQIGqr7lXz
jYklsrtlLg/Pqx7HzqXcpHrOX16aauFwD/fevKl8Ve7b0MstSoU8GnhJee7cv3Cof+bFI8TTi+EG
zearhO+KiSIJdp76f7RHLIvVNhV8ruTgbqwSscsyVhIXPSA8qvpJjssstAyYAm6g9UAJkkLRyEq2
ZEr8q6H5b3qfOPtEw0wW4tqI0dBCGckVgdk8bxhVGpZpWsh9Zyww19m13oZUjVZzQ2K/uUVoCwnC
1r4LVmZiBNSYkyF1aQ6DCYQcdYaUMP8mC5kW7EpByWn4/1ngj20Leb52rP2Ey1jn8028ZPBQybAw
OznbQ033S5VW1Fo2Eievxy9FRSqPiGgSoNf2lJk0PslOmc4eP6XYoC8MbC6Va6xGq79QlrgUQfog
ImVuCkhirSao6OAWK53znOydZXU0iDL9jS4eJyA6uNRsJQh197u2oUlOn9slygCKRHTqmjqnuw0D
fnt8onvBdY1W8zZorMHtcyRQDnREXFFt5kJNrfgELYbuX4Ru21oxrAkzyLoEgByIlYZhWmbQT2Ii
TfNUr+pWngEwk1/tdu1yvZ+2cpvC+LyM3h44RewFIZrbXhIjciAs+H8O8k4FC5HJzcS/RK2Qhu0N
ffPv7AGcB1Gpk5TdfkJHOIC+gc4c53OoWXZ6GOQdMQfSQHkTtFHE+JzUq3ENOassGBMJk6JzI1LR
pdOCOguEZHNx2emHTfb0HD0jL/fQ53+mAeylZxKIsjETchhcBMkkqBYUK86mlsdh8pRYYrx5M3Zx
7BSX/oFfKzAhbvCaQaMMcXfUYtzK5XYfjR5qyN9E1DU2uCxRTXuUowY2dPn8JMCQ2mh2Rh4JdLNJ
ZghV2Bs5HSjMjmvNNXvXiIhueSiwcogU+gBqRG8yqMhKLFi9Jgy0KqEO15/5XaDLQ2zsvnCYVyBy
GAVIEEuRYOqPHyPuJBErGwGvpk8S9mtKLOMN9na8rpar+mf2hkajjXRu5x9UUctrJIOuxdPuOVla
bcZDC6d4yAUNT9qaK6cYueqZug0hApMgO9u1ryoG8gVwPpBslobIQzYJEA2gvL90HiUD0CEqUYj2
eE1FKNobXcdcKtT9eIPLbjJkGm68w/TyVCAo/Hswnu4K8ev3nRMZ1yCqG9buSoqtLGPbdlNL17Fj
vC80/RVtiQhIOwoLiT6qm2vKaMLHM1yPACNq2dIYUihw0/gbWw8+XfFhAYkz4A7GS48nLFnntV1/
pyp8fLQHGY6HqKpI3WuSrhnkodF6IUaKwHcwij5MGxMkh3Yiy1MzaEYftj2+kJEeHkYKvTgn0s5X
/tBDX3cmUqfTtJW3PbiJb8QYxSuBr2XyOhPNXuiftJkpgWDa0oWmWpGhFGYaZJvv8roL+Fx07AUf
5RkqsTruTivdIUCzdAk4nax7sjzp2lzE/L10nYfJLmMWNMbvpFhoKVYhNyA3nqzDcLM1+Jsj4jaL
N9vapLDsgO803CYUjfma65SsrJX0LNmxTMOI8IHyyRr6CKsk3A6k1Qkw06cJaDTXU+YIa2TjiVEW
Typh2gTsbLPaTOnqYF1G9yK9tuqYuWKEMr1egwyShCgVHmI4mLuBV9fYk9tWERC9IuOC88jx9Smb
BB0kNmMmN8RSjAODOrGG7RiIKlwnXVD4166xNxwjGg5izzLIghCIRAjgwmbuCksB4Lw/iieOAvsW
khy623lXrvMrioKGBgSCe3Ra64j3SKlPeAFeufFUM+zYxIN8s3wzh9NveIwf5bgYhHLAATGozfE/
gWV06KsaWDcMJmbll/tqs1y1tKRWUGSfzFbiFdF3+Ybsrcvp7KY30+gYhqoCzKjrY5Bh3xloDG0n
4niL/5JXyPZhOUxsM57rvyYoUIFS8D8aiyWEil4vkNK4Esa1Gis//gFYfVhGR0eambBG+YVPQ9Yx
WQb3ogPaCPbB6Dbh5uohGWV/C3rz5OQQ6Nh8lLwQTftY6wJXaqY3biEzUKaM0cyGZvzuthG/Cztp
4HlKhYdcKQhHINiYEwBYFxLSOak7v6RPkvc3jy9hN7ScfG3hrUJg86W08b+l3UBReRmu3WV14G0r
yBf6tZ85ui4A6AtzP1Uq2geoHhEHLYyCSDePp/srLD3MNRgF2wVGWIJ+eyzCw4yUtxVjE8Jl+fxg
Nu89FrvrYQHcJCjqby2XbhSELwkf46MDJaD5RbUmqlpPQoJlSPycJCWGw3vlkxaNACWN73fWGCPT
RJjOZIcPGKD7OiJCMcO69pfr5vP7ouU1fW7IRh3ulOiGCZzXIIWyFrhfmTxgAiI/f/073rmiYbqK
C7kdJhBRMSjfEkd0+q1KOI5Pq7o56EVn+vr//W8crcvfLuDOy+nzXQ4mbgifZPBZIGgVx0+ujvNE
ypX7Ev+N6i9LON9GzJIYmXNGGB6l/nWeiecX/TFATy5BA4w7ITS1JbGAUY40+6afDCXbUliJJWJV
lR2Nyoxuvlswom2jHjQRLZnmFbr00YR85Cbg5iAOC9u0YzAILbhRDjf1wv5owaC2xXCMBskK2tkN
fexwAKRmYNxpEJLgoUKwKuF64gtw5mOAypXNa77W+tpsDTMBP3Akx867zOMIahHFa0JYwhmPvtvn
SuF/V5gHa/PLWdzUD887c9mtts/hA+yayqZfH1RMvmtmxPrIqw7vWB6whRahKZqSOoPsRvZuOizt
L6WnipPCbrYtwMNDMng3MJt/YCrBOyyGw7v/4OBwEP9UZXZN0UH8VZYesgdTYCGliRCXwRDaUXIG
eZKTj8mgMApL+BD8/gBuF2DTvYTgx8wYRrTgp1Si/kdD0HMHkawk9XIppeX8q9AOlVFTMh3fAc74
7+3rKPOGaFzwz2iVctEO08eYHDG/9h9SltdNeEPCxO6wwvIHasSOZ/bg+htVaouzCTFxjTRpgOKj
6iH7J59CldiR8qw7jMvGOvzXz5ZIOXqfkkSApIPfeQF0UMyFNRpC3c3sV0bCNPpQOUwTtSs7gUPi
JiCyeRo/X0hdmOSPfkDbTQcJreC/v0HTMM4M0KRGFhwtJJ1Wx0k2qoDVI+mIi4/tq16tCzyE5+Ra
R5VAL5IrKquUqvQg6yS/gqV0xwbG41rzI7ioWsdDFojrcN5q2xg4AjABt7p89yaQZi2XcaRBszMj
n14w651OE9ha1KbnKyx2C6DSV1JVXA3cOBuYHLXLvzWkqqlK+8Hsi6YZAlPWlWOdwWcn4m1Jb5qc
IS+m+LXcdJgyYuoJwwZw0Un37BQ+rI8S2r674tmHPKcsyWnjbPXFrkQoV/PPbZWuwnLlstEimBH8
vThKDLcSI6YfU+3YaQOEedr+XRqZDoO/5+FSSggj+tNDQdXZs0/oEQhwTJYNxs6/XR1ketccwgiP
38MyRkwG0KJcq/8zW3rgs6m6EHj6wpwt35eXugYzt3uRmGN3JBGwEGRf/BUCnfR2Uq9CM8WzslJN
KyyLpnasySwZKLWmQ//gHSGS4zDSAEMHUigSnYeZo3IYVWsTU5ZxRRRzdv0HGkgzPDvW57zkm5MI
g6rioUYqqy0G2cwpyVOMlfgw0E35f+5q2/uRcCEakrHU7wMW7OUwDOt8R8w8dcSNV7uvkbeAPf0f
IpnsFQTtxtYND7VMzdQMSRTGAincinAMLiYF9JkzbDLOET+wpxH+vfruyph1q1+IaIqeivjkk15P
nkXnKMUcFbCJpqoMt/XXlI+KywdlIqUo52IQITww5ms4bdq9gemUyAjzo0xPDGvFShNWo+OjjWaG
14l9PF2cW6TBanfOVhIi+K8r7IwlQtf/lw/d8Azc51fBY2bVGY+mrxYrwpsJbPxArVySajw/g1Jg
6ZVkb1YjRvTV8sTjeLvsdR57BnszaK/CoPOKtMEp8wD8dr0CM8bNzr5Rp206o1UVmB/HYTVbBpZe
qWRATT2MHQoC/Y3Lr/jX0A5PzITYVF4Fy/Q4WLC/AjRNJLa+U6xmv6w9bgHEishy3Pfi8aqOdxyx
BE7x+CmiH8nfdQsSH8aQYQbR5vGmgSJzZRv1Bi9gOupdKc1WVvVsVdBCe2SAMazESwMa1qkPg2BN
NkVllg8E7pwF7E6qyxOpCFXjdVJwKFESaAyfRE2B/HNkqwpJoU1VSnJ1M4UN3wDnfO95gNPJ8rAh
nMed7bZhR10lsiA3zvkdbc55oXqrRBOhYZOSckErOTLqO2f+4d1ovMnH26ANSNubsvUgikaDQmSg
ic0R9aQtXAWuIirhKodoKoynmKImHOOng4yxzTf0MidjEQt/b/Qx7ZnEy3VKrWW5xm13HMlY/8+x
sS7O54I8E59qN9gZtddxxap+NunNtMCKM+8wf8Y2aA07zPLLn+n1jj30F0v7y1hawlNMVM6WBUkW
MsxuzNjyBmoQf9SHj9oysfHBvKKo0F7LYUyihYNjtUcDA1y3BixIupSF5SxqrmaOjuSrGKeeV8wp
oXLxDW+72y+1X9e+uYoc5EYhvz5Bus5OvoCgXKDU6J1v8VWGX5ILyLLXEMnGGN/73EhCt05ZHyQd
XrV2a0/CKqWmEcwaPZNHcW32r4DMJNc2+ZXVUg3cF6NTirteTOWCegogeWVueLjlUNkCkAE3rV3/
P+gJ4uz4UkbPaygIYZixHOV6i0ZknbJ3wWq0GsJsdFx+3U8hMY51IGqMcYBpRfygCRf7AWArZrSu
NvJXRbSh2SycFiEUt3k58Y8gnVDvu7mFH9ZaT0KrigEzNT4Xr9VTjzThsNByN3Iqu7R4koeAibjg
/N06Wym0shz1aW4Y4U62SySIec4Yc5N9XKGD0H8SueVzwHQ1jBIIlekXesgrDDuEyD6fOp9UNWRW
6UNAAfUUybH/lOQcb9nuNsUnSqK4OFcFsQehSji6Hz4cxpil4zSk0YlvBjpFr0m4S3enS9RzzIsp
H+caB8TcXPgknCsJ/V7AGAFNJFgAUIVs9is72zchqlybQDUNKFFlezO3FT90miyK1+Jkt7moOniJ
1MrYe9YdenQtp19CX/kMiMNswKEpGr1OaIMaZ5UN5T0mQGRS2nctCX7sGqXkCQVMOXOhImA0Ym2W
Xb+QuFa9KewdC8ej2TYNrV5AQUlGXtUiZszOwzLEXQlZR4FkxKvVRmS7GLnCJ3i93WxHNKam7erw
OrIrbAR0w8cWTvGXynvS38ROTQ6Nc5UYSmQRF/OlaIhZDjkGXewhMDyPvhygI/sA68DXmg/LWYaU
Soz2tHV/uxDl9dPg+w5TUNMoC7/vL4tZEX7R8x7saIc3QeiqoXeD+dPXmhMYUlpl557kyZmyq++p
NHY7dJ5HFnmcSGAbxAYvME7M06iBhrX72EOn5ppaRmy2OvSo7vdYbwX2oUvZjsVVplsfFrv7rrFh
Sa5pNjF4jDoIcFAnmRqSARRURHxQcbbxiWyt22UbnvZOHGdfIqmh2n/YXKhFZX8OAMowiTmZkRLi
OpPRKVT5wvHYwwCzg3QU6NoOOd8WhIVGsXqjzfaGBdHHxdra+LoRA6J1cHiA7i3pq86lLNRwF8oz
kDfNMesTbJMBe+c5Wi7ZIfnwFz7oSBh3Tc7QLTZiVDSOzQF/hpHx4uCJknoNFiI61MahMH/erdeE
oMSJsaLDkbV0eaEYbTNdK+FWhvcqrWxiu7fCfLhVYSTZKz4coOdXs+VEifxEiCmichMjO4hRU9aT
YxOqGo+SDNauHdFK8D+U4Xbpwg4P+F1TjJQiQVpWt2kNq8UhovdgybJPbcJVvxBBKyk6KdCz51V7
l8P8826RClUDtWrOpeHogtqz8e7wO/xPDaMZcX2ZhqrDlGS1PzrH5b5VAcqb1k7MfJf17sYYSWAn
ctrpviLNuLM1uAbCfZayv/Rb5/bCLAfAYYjmyTSlfPU5UI2R4mbMuxdhuKc9h9URK2FmENipdRmv
kCDnydncyrABtPKH3EqwPABUbhRP98HZbfZL7F2pDuBNgN8JVPOvbUd4XObP6AYMXnSX6wEeaE58
pD4AD8qJ1ksK4EqKrqD+DM+8xIgwreDTQV1EhWFxkBP5IXXRHyn7okSfsXLNhfNWkZAnFXAL4ILG
D/9z0+ExPjqUNOwW6VNpcdQLXowZcVBkDYTHPugbxdiDM/o6ooEYe2IpAAC+AHtSOF3LpAc11adG
Ttq3Q023QzlFPD0Y+lJ0ko9jLKqirXvI54x3T6o2ELBG8TbWIM73DBIWwONvo7pd1mAoMWBR5wvT
Y/6Gr+Avdkpy3ek5WaM0pgL0WEesxxaSj22DeQDLEtbnRqKpttKwGgs4BTfcfOeERg9AyNEb1tEC
qxyB6FdYPBYAN6WeKBEag9uVS7xKL8UMbv+qmoheeaMd5G0iNbEGQ3BvBjZ86EmxtNIghAAcD9j0
2GtFUbCwXxo710Wknn48eCX/B5RA4M1ex2PfTmmMaFho9ndotTtFVJGdGUXswO/qHtzKj8CDH6Zl
zXeHh2fqMnDstVvUjIffS7zFLaRyXVGNvu7VwyF663YrDqRmtVTxGj93ABn/S1vKybRxpTfY7DOg
zVJ74BQx1Gi/4Ht9pWpbQEx3Wa8a24pv5/wrkYFnAstOhMlUDyVAhd0E430BxH0c+F8U/eRpAKCP
Ki73F5ftS0SYLDRoslHkBu70+zaKy/pIqPodgTFGjsqv+WIl6sI6ZPIMeQ83GCFXRywiEM9Q+osC
wGVwT1kzAS7bdL/l6vL97AAJy7GYhLH+GrrgPuxvP9yblCoJPbtiB9/hg/BUq78Io7YzqEMthauk
krjWLZ5P3JYgT9jy9sYcaEj6cnbV/abets4HxtgVFA8nN6kI2yVDHhx5IY1wgxKzJpFZe9bYsm4m
p2HIfv/OEg6BTwl5+JQR4z01QP3kdOboDpvJi84VP3ib4TA6EvC2iHaeE6nk4MCxrh02TW8txvm3
9Oq9TuMwHBuAM8AjYvxthxpkBpHDIH4yW2CwcMyPJXN+Ih+PUhF61hKPfxCTslOs/OsYO9SiVxxB
hAMIh75zSVZLkYUQAFWNMf8N5/+RX1BfAWuU5UjJQTAoXPcGvrxsyJ0VfTfIDIhfUS4Yz9e/KmiL
ghGNA4XS0i0SwLdHr3fhqAC+RAWF6XyR/jhx7hEvtS9SjhT2EDoYfXju/+RjFQXNcVMu96UXwn8e
JUlJ9ATZTS3lC8Hx116/17FmMMcr1MD/1nKP3cFw2lRKP7Lo5seM5zBszofjQXB0CA6xxNnWogCL
LObWaCdl/B5KPL/MlK/JQXwRJiDQ5bvraDzMvSXNB2vmhxmklcGxZrIasBUWDwnj19jx2SWs4Mr8
GJpSYUZfd65/ilI7rQdmRFMKjXdBjX3VNqiLiYKvmYMqYCd4XpfFKO0be0vq6tGSZFBbI2ByT5tb
VZRhc0pqS9TjxLUa6uYnYaHsFGTG+puCLpTYHV1Y4dbH3c5UWRvUDjHhyYeWbjl0DUZw57WJRpdL
gnSJxoZWlgwvqyvNwnwn7zT99l10XcFkUczX/KBawXpPkomGEzlPki4Jg4fg1HtO3yQrYhjQ6Hxt
2MsswFknmHfZp81HPob+lPILsZdOjUhYOHQfYuVFGdOm3ucIB098Gvd1ucqwpZBNQSuxOX+YPmKH
g8UKm2wa8dHh5wiB7yaH44/7xOHlrsjuNRlb1rAkluOJVD9uzBmTAe9hyMW1lwLJewAriGXLgxUv
8LV9kEn+45kB2tcOiOehNYHA4eOB614Cpo9kt2RZ3H0Mk+ApI/3xgLR3PU83uemrrrH748cpBwD2
xH5sAwXx0RgL046ZPp9vhdagma54B3aQa48jE4+bGAyKklRX07P/NZD0fJuWTN9owEsmZ/Td4ozI
3sBb6l3JLSyFiYajxL536mzL9BqWB5HgdY+QAYW6UWXvOTru8eBBExijTTc1WNMdPE93fEy1aUyu
dtKcpd1GcrOpAt57LIQiRsGxOdPllyvuPt50jJLMJzWagharcgD2SR3zsZVy5HoWPW3VvE8XkNWD
pSVM2PU23OMW3l9JTbb1Ba3YZSICjMR97jvts/fso5L6kmSahXUMQ7LAmtAbk8+iEsuuTsUQA7CN
J3cBopF0oDNiFx2K8QDht4Lp7qs/7DVgUAJXjoJgJ32Pj/B5WO6zUy4nJSsgmEKegYEDIRvr/v8X
4NK4P/q6wcQ6bnUn/J/Ss8ntcPVaUmJYtonmp46AjJNrOKMtVS36+67HcQa0wDQs1pTCIvJW+tCy
T412Y2AyF+nrWGK6YYiWRwSJviSGFSvoq+E2G1eEG96CIfBYe7kaEUu5vOlSWF7S02Y5YeSJOgJH
7lSQZhT46CHCA+Ff84tcZt165+3EHafSRNq8l5rJDDoTgPUNgWwlCAp1JhPE2GDc6elAx8wqAFFS
pmIYvoMqromTFLBEMHgHyxEC87Z5MO3FSbCNc2y9NIkEicbVkdRBYFN+X66SNgzu0y6bj8IzwOTa
0G5rMhspHaXLMWDhYTekZ0QK4JDj5k5divQUDoqODZhSxhNHgXGWAPwwYdrEs3P6Emtk/dxAIqpe
5n86bAmchfcv3p8aFmHhLX0LfvdMDm+0vZ9w/Ps5TcJbqCbLDp3/IGZ1IB59kVmVwvsXtJ7kkQA5
1N40x5pW9g5wJTSKfZZKZYcZGcADbLHnmqksvm7T36TEOEV7YIOdeehK5qmVGvpmpFvgG0ciJqJ9
x6iMRqHlZZzLyq4Ocza0x2jlwwzeYveQrSruM1EUnG+UdEj/Nenddtww0GdmeqUNZHYOwE9CBOf9
16tzrZLIAhrkZFHtfbAyGOe+oZii45GcjS2wr4/eAdbzWebGSKC49hbGWhh3Lq4qXmLsA80nd/qX
DeW4bZmcBgFmYvte9BVWwBNtkwz3c/8XcS1LWJM8uknVISL9DYD3VFpeqLGxSL+N5u0rs6g1/oF/
dJcdUPfprLrqevG1zAon1xfe/ixGMDaYj8X5y0MbVRakxMdbYr65UUwHRysW0FQB3A5GjB7cDAoE
Gk5r113PAqfJICJu4ddQOPPTP4CNG/VbhHb2qZYHYwIGQuqLuei2LpSHF1Dy3lXyMxIlqfHWIt7a
imyZUAoCSAMwvlItbik1spBvsYWBj8htwc+ZMcbDBHBQ/juO90ZdspnQF6EYTImCmtI3ZtrK3JP7
006KxDR7HAYtY9i1D0HeK87hj+69U+xjjPC/AUyBZf7FN8G1o5tNmtCaaHAgwRRHmGA+0tv8an4i
ADEG8Jso4pPJmEsxmvo7K4cfi2A1sJxmG+RJrVn0IhLLuqXaI89SsmilaaEOBQQRVEwDpUJA0Vzk
Lt7Fhvmp9KKHvq3ZMIjBJvL3+OHFJeumVJlz+BHbgsOImCHY8ecG6XnXqxsoKJTnHJshDyGBsXGa
/ffa9I3u2Dqb1JdnHVX5/8rZ15AHxY/XjDUFpihTMmw9yfw9+6KoWH5oTiRnlhZ/bI6a7jx7xGHd
zGdH0ZGiCT9cV++T9cEzPZZQZ0aEfYUa/1gc5yuoEHmYJznlX6FsCbbIcDMe6nI5KU6CzRCOtQRl
d4IXFJH3jDQjlGeBt9gzlpo6lh6G3fgrlgdi+YeY85RYczwm9PKtco+1+RzRbCNi3Gmr2nlgGhpR
v4j1qDTb940JmSENFwb35gq4qQgW+QnJPWomfOR2FrvkND5a52xKotNy1VfGGNv9Zwydb+sSwegO
FSTXjV9o7GGTr/cnq3mdFKxx6fQS03e5MZA+BIQK6RfXt8/FgnBBsKd2xntrkIFBN1AqVMX51WrE
H9EjlHgbVs4N8iwgGOZfttNq+EC2vFfio51v6KkBbVizJWfqDL+qhHIQFxPGHoiv8XInP/ddLZqg
hl1Obp+AzWfffTeW749V4X37uETfNeAXu8Sl+rq5LQ/x5BiQx/6EPTrhl1dLqpn3YO/F8fVXz1+y
pMY4izJvmSZX6A4gVmB+6i0kJuOr7+3SQGaW/w3ARHzqka+hVznoF34fekVnc38i7l4+lghApGlG
qpzPWnGA7NH/cfs9upUNKSPf70XqJlWtM943ySKciaY6eooYFaQTu8k0cOMJicZrfTIqV4KnayjW
xHGnKK5SlpyM2C42+j+6l0HDszIrgL9FPvv8lkA8kWX/mupXuxU5E7ZJugBL48wocupIfadSq54I
A6EmU9h7yGZU5bZBIhAVRp8m8k/tXsFlWGwbwcFOjMK/EnfUc6TU55t2z6q8pAgDd12kE9iCIRt6
5Ba9sTrlQttlz1AH6/vU7FPz9ZN/h2mVKubX/Vwik+EO5KUCtWq4eqfpDTfy7n6TxmK+bxI0Jelq
nvtW8K/kZScHV2TPW7Tu1g8rzr64ZrW7eu6M2e1FfSATiHAC3hk+0WJl7kiI/nJQnjjN/CRGdCCC
v8Y7jE6SHXB2CVDBlXnbItlfw/6T//tjHQTpceVlg+zCTw75YQdUEe3mk38WjpbYqpb8knCG76kL
fs2jWRTShKoU5zBPLkr9zbXqkd5W1PaWBkn3pJy0Eynjr7eP8wjvlv7QU8hna6oqceWwWcoSz3SL
5BQdXx9ZvSjYPMaKFZyLbjnWS4fDt6sjVPeOZ2ct8uEcJcLn65xnlMWSgbnSHDVJvVDuCkcs7IbS
9F5YZYUOElkP6O2n4VBtB6EoBZ/mM8GgpgGuHSKEh69YYRXSOnOqGe0UpKLFLvAgK6/KCQ7UtzV3
bRrnquCMtL5psUapPGp0XSzTgF7NCtWq5LSGFmacvDOGsv+9Pv4mzA4BDo74dkZHJC8EUZlq4jUh
gbWN7NMxkTsDAzczFiZkoa017+3Jb4lil1qJz4lhSIx+343g9X5mHqzM+6quXf5g/JG7RTNq5uKK
02dyqW9UyI9zPWMnZBFprSXBo/1U7DEmrq16nvIABlHzN90oMFKtc+ByWEeK7+12Amfb3Ws+LJDX
vygXDXx2oBjx5qt8rh+99y0dvkJm271Q+1fJa5aW4ZVPSE1ae+xR+h5VkRQKP8ORdo5kW7Ayseep
Ddugaoy8shE+RaJKXoOBbU77Si0Dpfsl7zAFvh77MomiLbGGOMzuid158Y1JzGtPGuY38BbUHdiI
fyYSxHKhUD3XfO/Wt5gcwaZKdDOUaFxkjMk7/OhN+AJxvUa8ZYlIM/IDtj6RFXkpYzA/BLB47su7
lXGQWZP9kT7ymDeu6o3Bttzn711BTiMf+uHKurFTYMZ7/9t+9rSSMGobl54ClzgrhYToPyTEYXA8
mQCqIcIs5Hn3cdybeJD2sD7QHFttZuKxrQ9RSwpRv/bzHmubSSiqlTq++cZLfHR+ik+0N8XcoEZ1
0w4Q0bsqhmUp5RRKSTqj2aZVsk2261hDabO5bUx434/rruiuXTv/ZvbGSRSMipF/xmDduxIj0UZF
SXeBPplnon97pq7TOihMjVGMmr1oMqxCemI9BHL+b2PMRLkSPepQ9p2IOjVpItfkssgIkP/Mk5qg
64iEnOvnMmpO6hMy3Ic3o47hsHUzFH7HvYvIcK0vj1LC/Yv/8NUQ2vSTQ4NJS2HNv7zMaDA2GUHi
vgqm2rWh+Q3AGgb289gUcJYbnIPxR7+YR5DMxNdVhPdLjQjn9gnU3B0+CtO1MllZ3sXXdX6lHLaV
dpvhG72pluPwOgH8x1oaqyWjw5ynbUP9dBeoM4+HiPM06h5GVkjVm33+dIJ706pt8s2i14hlbQyW
3cyB+vuZnxaf4fDvJFbgfsSQOwI3VrHkhPkQp6jvnVm034uoO6qfRosFM15R17734vrsZbg2USh7
WSxZhoCgeDONg5WHG3B9YioW4++WNQBV+YeLCYACubpUmTMNjQlxG4nfrOiN2FUcPJiKRTED0OsI
wjbRL2ILUfngFcLWMFbds3k0OCiOaQU8OPkMwDKy24sEeTkIAazmTCHp6QOoYvXpQ9qpmDJrTWcD
m0bSlQmhTHucB8VrQL9jua0gNGt/22bVUrG7LSAWdbSf02HBe3/zPmGJbz360RrmjblHIk4YnrtY
vfxKj8+9Ah1hdgnea4xxxjkEIUFmygaBvs7Yb7I6X45NDAe92HwDadzj3nTvgn6WPQBMKyVH9Mt1
n7D/JMd+4Ef3Iogjlcc08nF3vue7+a5A02FIbtWeyIKsy/5WUEmyOS/Etn9tOqxXz9Z5aj/GJRDP
fh/xWyZKz3BnAzrl+8mYgNBDOxLD3iEYdcnD4Q1SrUXhSV0Vx6XZBcoOzbAXQCs8nK9Us35R/i8I
/KDCAa54ajFMr20ua5Ibb9xvf1C+wHjTSmHBKCalsKqa6td1f3gi6QHz8U2NAvka5+UzgRxUOzo8
C/hzEkGjW3TAAdqFh2qcH2Rqr8LcpUZ9/71IkNoD8qvNcqXQYE2GIfr2MZVjmt+nYfF25MfQjuEl
it5Di7HEfx1QyJwVRNRBhvTmB70Ov6hGBou8e7Vifrx4vb5stu4/51s3elZs/8VQIfTnx7lvLhix
Yi2B501By9ONoJkDtDNNmGuHaBcikwqWKEWhVCQh9HQqZMjzevgHxIE5eiT9u8ZTBXpc3zUBjOWW
8cNgdFXBAfDN+TjDCfn+FY4oY/fzOakNb4/ozgznRbImir2qcDnM/zQt1sFJh2BJ25Y2Zb+Z8RBJ
Y85HrxrQzHw9y/06SZbYSEgwiMpXjgzJg94gpC2GGjl4H3vWu5b+kcsKgdm8UTVMMT84e2hcp2mc
hbJfUjYFulAPmZKyt/AA9QKm6R1ZRx08Lupzkmj4uV7U6Pu5MuB4QlQ1IRfN0wprD3tDT1fokEQ3
EKVOL3NiJqh2JvWnLTyf5G04Iflc/L4QkKDkTh9EYVaoVqtJk713LDJsGVbHFbVYbtGKpJCPyb7q
Qfj64y6Gxhhjujtcj+3IJYCHmpL2Bz9b1na6HjjNRzJxfqIonkApkH3cKO2ZJVl/jovkdvwGv60I
Prnb1iAzgD/Po6YNBhktpv/cbdpbFWl3Ye2Q9LDZ10MSkteF+533oz8hORokqHf7Csp7AX7+t0Z3
x/Zrqv4P/WcbRmeqF8zumEqWw30SJPAY52A8ypqkCjkd6PBdk7PgVn1RFkCi8AGmpDxKSbC2uxE7
4JlU/mfsL2cnv+lJM0ubM4CN6qo8hZ8sWWDvK5IbE9kooKAnmyt1aPXd5HRn0ZEOsnN+c2+9rXWq
5qvGKHS7BI27fA1uGTwDTiEvYmOkQNV50gg7DGa8Ndv9+Vi/iOFNNfY5UgbJO4h7sil3OUJTHy25
gmIlVMPDIOyRGA6AtTYXF8NLiQ2t1JHZcCBDzU9xzL3coqxA3NHHegxxaL9J/MEe/1/J3LN50j/p
NdiE4FhDvgjcmx73a4sRrgzicYTU82iSLOuwUPaxRIxQyjoA5E7m2lTNb2M+esJBUgQHDbXIDpL9
0fcroSzF/7g/hWYxGuWOnXPMWecykUhkY+N5A76ondNN8MtaX7FBoTfRaEv7mYfgMFleYofgI2oA
sm1nMSTsXV7C7McO3bCV1Wz1LrfxRdNYmE+z7ChtIwd81gXddLiqD/jn6oSl/oHOl0SpE1flde6d
GqDtdMd0PckwDNsQT04ekT7U4S3kQkpyIdn42tSRrlEcY2IykoA2S/pi1NH/KXOQqXF9xPXl1Md/
cc32jKZb+q44ioHoly2DJWgn4LF5INlKprJpVbY0wSOUFu47sFwtplXwUHev2QIQOiX2cyAtlegD
9JX9gWwBtnRu0wZWdMBZMifo0jaRK1ywxi12iyzAihmg2yj77CZIeHx/7HlEvOU7KRieq220jonV
EQ3kUqu1RaQebCDxWZA6q35cyHAucVl7xxxnu+pv6gLsQudLfFR6+0WyM/JYxv23vxdGl4RabAot
obkxdA9nSGvmIpzmeVpFOECq8mZokE4KqhnAvV82ttk4b07Szw0RlRnhnnxx18tNFTBH+RDYLjmc
BncPXrskhf8EDct3rzRBi3/ql41EVwxPOGCO2pTNBMWEPjTSZ9qFNUktFXzrMS3Vhx+aKM/SyCta
awNkgURn0XHtGMRCZW/60yhWWVi+pVlRBIq1i0REWzCisRY0+tHVkcKs7EBp2T6nWjuVonpVZQm0
8ReNc/YC6k8S74yCJ5oliBZfhgwjK6fn1VJ6CcmCd2jJyVXtf4qcJnGKo6/aRqQHOHd10NrhajN2
Su5KzGWj0Z5XYkfSMpAaac/phfV7Ngq0mpXHHWfMe+jIwpqTUJXuzgccfv/0m0+dhS01uARBi0Jy
P+0RO+6CxpC1Tm1AzL/AH3LBPqHX/vqs7uYWSWvFye1lDorIq5O47xdeNvNYnL9FwCLETDE9ILSb
a10bqRvOPZ+x0Y8wQaZpmowjizJa+4QebgwRd645ZwUo9gus/pZpEqsBcyjlt2jpQbU7r9v+n8xb
D1oGcaiWdt+fFQEG1+AryZ58nHGUC72lw3bPKcozCz1+vmvEBltBXgCIB5UOviQbzG6omzGxntX2
uzwWv5n+zlTI4rKYQhL0swp4e3zIMxdAgYMHdqI9R3a3GWMZzix4+9ifcgoanGmlRvshSPKtQ+ah
o4OW73IjJSeVr5h7ldxPH1+lquYyiXtqxMIwbLqvEiBL4PLV3bC5dfUGVx8eMLTP+zBGkdUYz36b
pQEejUU0glmiIkS2LjmfSonTZH7zOueBBCB6JpGe6BCLJmcf6x4Z7+Rr1fp3wu7Mz9ZHg86HdlWs
vLr9iMAl+MtzPcrXybRilH4BbSOw5x7rKO4rvAGEew1hRcPO2ODrHjgw97DD9PJTX0PFrciydsn/
yeOTBumOdQxzHMQdgjqHunzezXjmpLyAi1+awv4/g2h8Dbkt6fRxjJEixX2toWRHnA/MRhczo+J7
obeUuM/kHsYhFMrM6009ln9aLesMqI4fTG17Ydodb/hmb5cs044bRZ1tuOnD143sUEA7g5//z8Ta
Zw3+k+9goY34fv1/zPEbA/Nd/01gyBb5dWRR+2fvs2dru89nlKdgmj9CLaBjNnX8hQv47MwmGisg
20yzIrqOUn/jp3a6Hom6BewCklSY1/R9zWzDFyndg24Pzgm/Qzdh3pNGl+smcR5OTPIIFQEFGKAu
5o3dHbyXulLKC9vFxg9LwkHGj+hIM8yzuOIzSfcmZT/BJjq4JQ8MmgpAuXDx1Ad9402wBIso6f2Z
9/8Y1AhXJSh1ZSUMZa+npMmpzDTyQ1kQJe9shXQ8W8YpvVYCpgY/o6FWVUqXm5gW+P4bTeFBdS4O
dFHtIeXP8O709ghAStX+wEE72YxYh19+/IzaLjgLhbU3wjLok+0+uk9bwhEypKxmo/L86kMcfg9m
v59mQD8LQS9ZrkibuL+HC6exqqKpK6hzEiMT4JaChbB3ZF+m0k7UxYOUXGUYmhLGbJp8EcAAn6TK
LzwJ+4fttMH6cn5zk03t45tx2dD5sYGvu1v8FYuvWgvgbT5iO3aYztMfKxq6yuKiaKfeL3T9hADy
6/st0IdAW1AfMyXEG2ObDSvZplRfLsfvafaSEudkNxnPR/whZ1ihW0cNol3hZCJtdJ1ynJmu7r/k
mqRL0LONsdph34zBB7XgyZFSZjLy7b9rln5PDC5nWxuUz9/YlSu9/KKpU/HpF332DvFJMnrzwB9x
NsjbEPaqzKhMIPW/XX0LeFD7IfUFN8WxykxAICyj7anjCqfU41Ov5Y7AfCXecUdcdikKX91CPxgM
mMz7XUdHDozIblL7EnYTnGGjg6CgHpkPwMgIX2N1vh7nHMVdJYCpppZ93WVr7FF9RduTft8acAIG
RxyzjyjglgQUQOpS9yecoiYYBDQFHlu0Hp0413R1ruoke/nevbFFdNtkkk9WiFfTQSOx0DwJm5lL
CvQagimB1QANj09HoXycwi3fL4s2hrqsHRl1L8xsR0ykdlgTMjPoyVghGtfzrdkau3OtyZ5mZ6Lg
ZFn715KXAg/lromdFF8byhm5nI7nf9ASTOyqgAX2KaVCuCOAthVpJhCraD+zrthOK3s9TPAjqW+g
ZCra2ZeP+wGniLX2QUVbWhrEFg0zJeStFu6UoOve1F3Rk5ABMuFRyEuNSek6Gt3ugm1251VNy5hC
vweDeUKdtJ1PBKYRz8l43nPOCqAryFe2jVC/AQY2CVhe5dQCQZjlpF4ZqV6yDPwtKnetGoln8Lpb
oQ2Xx6kzwcSiQjqto7Dsky5F9H+56Mz5hE5C3ketp2KlI4A9RSuFT75b1waCOYD+XzU0eMM0Dcah
5xAona6pbrwQoHXgseKq9KbHRtZLyhxvea4I4Nm8lgzwCDkQd5tylJmoIY0r0g3bW/2cjxbUVGUy
P06iFcZd47IJOoLind4OaY86HAbMSCvm0659OaSNZiAIzScP07Yj74bF392ZoCtbVh4GUzDc8SKZ
u2rzb9XhLhY/2tXUA6Ujxo1NsJ+tEms1germ/z0fRotfWfP2YmRZFR865ETJlhUyGXh8y6E1sbhF
BQEEM2xW/JJXMzvNt+FlMiSIPw07DiYXKZrVn4FgqBwXQOotA/ugEkY/B3JDiNR2x5vlQTKeD0Rv
o2jLnIgCX3ocM8iyeUlvoCFQjB5A7eOJazR/RRbiVdmhqGlScZLwu9MD8rqXOKh1NluySGFHkrVN
5HqSJ3XucSaC2Eki77GrN9hjYOV5URlOLq7YzSK33WD9e4ZXRg5HE/DR/YyJGZWGk8ZkLCfhd1Mf
XO2hhAFX0pHJavGes9uMJ8uv2K4WQJYnZnBRYKYG8bA2QrLZuOwyk7DHlEyjNw6erLnCgTn4KgCp
Sk1/mAKyuYa2DW+0HhiKmgVLuDIpikZQr9XQNiTMkStx1knqLW1t6otDIA4T5h4qoNUjCc26taue
XizlSKFq0OsNz5WvvwuNHVmtMynKTliRQ9/PD4xxu9pxn4C0851ZJXMMZ6MEhiyScbMiFWCQqj0h
IuslX/zEMWNPXtgPayNc6S9FerVZ8oM7GsH7mB8uQNYY4mqzHaIxGIbV4EqpoJcZDPib1FQe4eRG
bJFlbyshuZZkqSh6EUeyRw1OP1OA7MGbNsTsHAwAjpnfliGz/mtAcGO8tVDYKJj4gAAJObPkemC/
4JTxh7nWRi7pUmOORE+x/kWSvegEoH7MN87QIrcXVOyTJg03uI0GKKv8QNAdRQRYQXz6y/sb/EGv
eKeXsVh/GfHwFnCLxnM1w7GQL2Vy044Tattl1wuLrJlfZKrVrKp8+APzBJibacokMYZDsOAgu/l8
AgKE+lhKxCPNTJfPDI5FA8XfUs6BotOm9R9V6d4/bl380CLxHYzzOPgCRh7wH04Sb1/aqkcuHbJf
pgSrmyKWBDqzLof9J02ba9CiM51v6LjPHs/Yg1v9NmvbprP3jBKw+JwxG9Dj6eMQdWZlNL8VRA5J
+7zd8dher9+R/VRB5BSSsUqgpi33tnbSvtWcyDz5PXeJUV4IgMfuPYc+amOCzMRGaltt/RxLDrIQ
Cn9yeXSd+gNoinMR0TH3q4cMhtnHMIJZvs8hC0OQfCx9uSUH2HGzWZ4k965GpU89zSibU0iwbvWx
pbt7wxzATScEfFxUW7Ld1E0hcpJ2dMl57e9SeRGXvw4FdrQSxNr3PhwBgWwGBfhTtYCCiqmgA3T5
EbB1J2BcmmqskmUskRwNiI+OzLf8ckfdfBsyWJGGBBdK/OB9qkjQ8zGFO/qtxBNaulMNkA/aVtA0
UVQGo3OkDhYKbPXm12TNaCOoeN6DHENiMzuZSaik30NQ2anAzuMDGeu6rMzz2TMWcmWvCI8M9s4c
85rSYOewIecTLyB3X/DjtHkSdNkkY2EvF8mlIJuhby43UYFVAO0fj/gwU6AvcoRcfkI+9gxqzyy/
4TwWRJfIvVVoeOVN54NuVe8qxZngivJ/NhlqTU7RYNola7TkJVTZXORxZSEZZN2xvD/BDI6uI3/R
CJvCgXfbhyqwf/QbDIaxCB4TFu7zOdZbwoLTyUjgvZc9mCTUE8PNbv/+kLZpythDAJhMup4lmDUR
g9Gs0c08FAlxLm55ECixfC2Qe9PTgCol3VLXW38MX2t3oEuMeMKv6tlH49spn2ROaYL2tqLD/12L
auBHciSFT7IFwLXHKcpnM76bwVUN0+dxdQjRL6E8RH73d4/jTStAV6/2OMLSvmmN/QmvkmTPXUYe
8z5VGOutlVoZdzT1o1N4azR9qZxbFmLNpHfc0ziSRLfD5J4OmJEgmsYB0JAe2cA9rK2GZ8dwb06N
3NUPj0BHRBFAtIrP+gZX4wi8ep8qIs+/JVAedshDF+qpcSqQp1fOoUuI67zRqL3UjCrX9BorBTi7
cXH+jqlzKJ59FLttp39ywIx/cIr8lSQa3FvL6s7NaWT3DfPcgAj+dmrAsmRI9gh8jKOGCjaaHj5j
+r/ssk2Hm/YZ+t9CakZdMKNAoPDs4yg28RImmdnrkd1hKkHp+Gvm1gcsEJEgguf3Im4zo6zDWLVs
t0eUZ8CzebMFAPgiiZUEAp3FLR0dPxRj+8G7jcDi7Ik6FCSgIrJAVOf+K0q+pcOcoXY+aa48U1qJ
TePV/veYZRwLfMxyxqnFFCJyn5DKJ+tkBMxD+6PXMFSZ1vM86Elpp3MbP/Y0lK35W3J1F9WikBcR
6G8RobXlRkz5SE0kTevNi0cAvPzAEABcWzvexnGLObe2Aot8/2pXYTqSJhS5MNVEJ9aji+BjchZY
BuJbABr50kKFtBgOfK4mncJdsK5RM5JIEUBIkYzm7hiDTEv0Nx85vsmHHsvq3CfmY/XX4wy0cNZx
k6BUFQPTMnsrea1KaJKDDaXq3lPWc7GIbYj7Vb9adWjnOc2xRO3QLp0708WDR72LS9dQGag3prfS
l7OK1IDE4w4yqyyhTD4pNhXuAcva3mNQRUAc+A3QZpUHIww0+WepzMgCW7gNuGsgda3F+SDPPIol
6QE00UuddnpfV7kuBjkNQST+Naf/0w7KDOO3txO4QfnD18b7mhS67InOIr3TYmjCkAde93MB52gr
4M1eqZF8ddjWud1oBv9hNVBpwKOpKPyfVq+IkSonpCZEWuSawI8NOo5NP8Jfcjk/tw4tldMlfSxk
g8+twpGvc8YcavXAXTgBdvG4mU0dZQZ5LCSleLAiLB2Roy6NSpxNC1O1aSom973e4TPApZEoY1iQ
EBc42mK5KUNCD1+Nm2DKnmX0osffImdiJUL10T1tLxtRSkz9avflQrRbr/oo5XFX2y6wIbgXmyk7
Oy4onZQjW8g9F97+YYXhddaqBE+vk4g6ivtTJwog1tReMuMe84EX5jXdqswx/mFhBnnTjsMXCiyJ
T6FePr59m68/5WJGPKVDWPszP2pRt3sajSS/Ywtw1C0HGjD/XIcb2JfLfTLmh6lPk3vVyejVIvfj
nv3gNHYtULQK4MODweA9u2p5Lb0YYMKd7tVv3ZKEzSnlyA+mJz/srrXnz0mEkq0DWSGd6PeDn51r
+UcsXp6Bh+iffuoKs+3eFiusQtJDRapIxyiAf8mPV3UaHZV6zKd0wmIWTz4D+ajNWeJ+7QOmbkVu
OiQ7TOf4NdM4ZI1T+e4dTUbYh46/pi0xNtUlxu+3SHIBc32BAybi9Uq4mljYcnJFzbwCOGsp6RJb
SJUwaLGx0z8VuOEAJu2fdaybE7eoMFYcWRe3RIRPkkQh3GUO7lLhWYDPSLSAaAemsEM+DJzG+InQ
Ie7ufavH4m+BvmxZL9HbB0sv7Rq6nXpf0B8nV9ESDFYVEedqKIVuTBWMcO1vcFDoB5O893NRfXzL
MrE6lFI7hzZuc1LyX5nuP9AxP3g4qtjEiBruxfJBJ9A26gEsuRVQ+kF5wggYhyP23876sO7bChSt
S6nXCOSxTYrqrXMFhDYdBkz3GbxR0EjeZmk/0Y2JR0HM9EffWyDk7RwerSBhr3GXtqbMyb1QEP1H
IHblGBjR0OaZVXv9/HIFFucWkezIPSH5qbeCqnekkbeISkRzBaooXnkS2kuLxkiGkNO+H4IPEQe4
q/ZEVqTpjkvRNc2Xi1sjZGxPK9NRi0Yv3L7neOuEzk/mJYvRwmUMH7hxIlM6RiLEByvrYImnclKe
1+VRpA4hSe5pv5plTlknUYUoK8xMgnQwn8bjalZjOJtyiP3uqa3GZp8C+e2XRxbkK92GZ15jkHR3
+S/EbtDlBZxnQQOjXtJji/92tWlo0GuZXxQl7f5wl/AdfOTOYX9OMhF8x835S43F/017w/zbveC8
BJcf4T1pchZgCaUcyTUjcWjE346/V2Uph0R7SmltizK+H+fMaZN5FIlXE1G3JNX/zJ6JeaCPwfCa
mgriYTkjrHDse/3kht3H9bYi1atcqPZJtZCGCRspN7Wtw5HRLho4JpbD39awCi6ls4V4yDkgm7rD
Qwxm9lac1vZ1yy19m8v8+NUVpSFCguSBcjR1QLL0ouH9szPZWHHreH9txwKxo2zjvKkrVX32oLFE
q/T+r+aDefJP94IyX3pTu9iDT05IiNSS5ERPBxYWvgry6OlUbmEAukMArPaGRQZO6muauRcJ9OH3
hqsmT+P0OtqnO4GqT2Xsg7qKbcPg+gqSOBxLc07UEi41OGP2BkMZ4phNODkCkyoKv1MrzhG4yj24
er1z/yX0mFXvrin8mQQ6fc9ub6uykXpZUJcmbGqUDlSYnWRkZv345pGKxABldaSpxu+LQCKsGaJP
O/Wy2eUzN0kxNWTNDr0qowyldHoESvHqmpK1DHWMvSsCrKQFsBCezyNx3fpRWPyXtkbtV4UQxR5t
6XNoLirAXTdtbaBmlPGdFey9WtB6kh+5BGvhbGzAPF/zNzwe45M2lvTlL03ylGWV5CrOJvgBh/gh
2p78G9hHTiWb8QUuMrDBe/6un8vHUIzk33Z6zga5iRCV9snXfo+Rw+P8EFtDSBb9lvJ4g1g8BME1
PkyB6NORsspPXGovwQ39MA191eB/eWs0uS1X/ms0is68lB+mhuXcYdYbgDFVrx7pNLRKgzI9P6v1
UVKl9l/lH/FNRA2f4DMv4/SzZesFM6cNHSib0d5PK9P7JqdA1MImf541SH9e0wG/SCUMhayLTrUo
HxRARlsWo28UbJyAutf2f5nym8qStx99PgmbdksaqnmHTo8hUtHrYShOcH7PAK3JR87LusrK5OwQ
bmHRO5i4bvwDFKAD8vtTDVp6wPhjdz4OsH6VWvNOZYf/7DKPenGjZv8Lsd0S0P8GMNge5P30jCnM
kxkS+5Tu4TAprcfckG0VS2xej68iQ72QoNjCfx1fmPoeye/fcWRZprZpw8aAtvZQJkKGAvw24UPr
vbwVUV9Wm1kLgFjf0udB9nkSfgj9jBTcJEFrBslgdpUYsu+bHkbP2qonDf6tNK+Tfi7UecuynQZX
qjrxDPfp/6NhuOyWnQhIEdsNJLevcOR8ZGaIwhnrP4RaXmP/ihlFH3S7rosi7gwEIYXaYQVbX2k2
2qEBDbPM6CKFrhsNl1wRP+ZkMsWkrMQqRzlbfL33pWC9LtN4jqF/79aPaHWHqjNZjkigEeEKe12x
/TdrVgve6f/PWCtaUHbnfbAT4rHbMJqDH1QTuzn4aR9fiaiVH6KB0NX5cFbmsXIqL4ObtGhSwYcO
FaTv7RZaoSNVY9ZGXUpAm7rFSPBK5pSLpRh6AHD0jHpVC5DSUTAxT97htS0h1pkD8kKBE+1dmg71
pw4cvag7QWV6Z03tS26GWoCzNApKMyYJMyvDFGZGDBR988iNtHtw0NeaRo3qwIGAUTuHOWRIQftL
PLVmIeDcvhCbtpv4K4XXqrhPHL2X/rUmoEwYMCHWo4p4C5ZHK5wRPddo9YsJjajWv7sPNrYB8cjk
LqBEfBhuuW2TEQRYgyHCNQTjTr2sTW0LuupfjpoF7qwwe1MioOtfyfINwynK8t64JUDQH0W+4xwZ
Xxq3Th2vDSyZ3DKtbF2s8sgxr60QU11huRguGrR/AENERWdf84XPowj0f5RJ1bADe3v+lH2N6jNE
UFpNEwWNhBamIp9j+HTPekaDCzjhDVzbl1G1D/ufecXv12tnMq+qTJl4QO5ZCIKTbBTWh4Jg53Ts
qCHYFc+Ke3XGg4TtIQITYMTRlOr+wgrD0ErRLLPCWwcHDHTaTeu4KyaIiY3BRsGyzXTfGLW8n+bN
H915vDAz9P2DtFAGzSN5tcMvs07N4BKsYjMSin18vqxU9RBOAh31oJ/SzSYT7Mq/17JB60omkDta
V33ZxujDKWMtRXmnxE3PvjXFMGmIrDzO0RbWUBPrgnlVN7fT2yyd4sxP6Ts/xY5qriL84pC//oNw
9Chtme4TuU7ZI1Tc7U5GQnzLfzLsV+tJvH4pKVb+dU6ofnyqPYAxsSrffm/NuCwIbkIp6yDwaZIt
a3DydsKGRnWtOcAgvOqZKg5f7a28GBtjbmDnIVYzEJZEPipMQo62F9J0Z1092zE8pFfmSIA6YEIB
lWJ/Tz0KAmvqHRKaO0g/96g6Pz4Rx/nMtozrHHfOQ62IdXW+mt6FzY41jIx+GaObdICppdCIe4uo
YDgEejA9faq0M8ADwLD2mjdZie1EsouMMqceT8zmkNa6K59B9tiEpIsTKI4RbBMP9HMTcZeE5qv5
nKjCu8vaisTTi1s9cxZlbh3imj9/BlnH65GZ6iqG6xvGyuwWLqAwufTTxDZR5BYl3Stg2uMi3oU4
6Vdi4U0hKI3wj4f4x1fAsZXTjFO6VWiHeYyb6IjpyL5sYiB1Us+aI5j6fRuV3eZTJADKLAq+EIFN
9gkTi0WsS12FlHbshqJKoC8fiGnonEghD5TxjAsXgm3ahz2sxYpvAJ2SmFz2ykRem1u2i4sHHcKM
3v0qW7rRXjYaMyfU58w36z9Z5WdOGO2TOidOskg7x4K9VodmMUICJXFnnaI9k9Y2apwEYa7nHXia
7zJ09ADIwW065fXhmeIIlj+FrbLgcGolt6OhrfhUliAZiS9BKoaodX0fF1Fiha2eBr0bWU1ixOzq
2OCN7kSu4zYTNS1CQOThVgNVo2eYWoST1Wb084IxJXGPBN4uulpBfs0NN2AfOhwiJICHg///O6gc
B/3ZbN4Jck2ESkPDCW/7zkglZQWqF48ep63gZAJEnyjiXYiHPl9TRg61q5p7GSq5U10TPy9Oc/K+
Q+GLZRpZgSEXyozhIFNdG1JQPM1Y9jsiODJHEaONeX1VQBz6RWqVZgLdPQ2wGcl6PVih20mEfbxV
rBq9rzO+ISXcufnKclhjqU0a7JFSaEH96cWWZW380398eeDHrdLRHhJtOMdPNQW4aavIyOvzdulc
cwukidXv7sxEsmvgU29zNOhGC3DJF0OIy9hM8pOnp/y32s3Rev2UQxhmTxzPDfADW36SEt21BvSv
95Zke4R5UJn9j7V/8dWNj60H/urKi3BK3ky/Kt2HLRH+48v2GpcVkZaEzHVzOBsaDYhALjYyForu
OKMN4roROsn7IbNbTyHz1bpo6EnZNOJmdjns6rcGGdU4Z5s6ZiWzMLwioCPiUZEykQlUhdKIa2VR
2Ui9WLPnBNAySrCKVLVDayom4tuY2FirxF8LyZvDamc3Fuxrb6r4NW6DZZ0dnYL4GsazS6vVkOBW
jX7QkZsLDiwouaB1wcrJxrn9bp23Yh20dNos3wurDqNQhY/9ja2yvJlJDrVNf6C+qef7F6wVLv/Q
vTkBNZeQ6U/amZpiSkYiStt0Cfeeayg/aqGA1XlsYXwgMPwoZYMrJww9jqw4Wbfmz3cLjQo2eERP
n5DdbXGyrfwn9yBLoTtsu1oWsxc4UmvPRwDzcQsoYNFU4Two+G4oD1TBJjmIgxBgHejNM/fzv+sT
cjNgtjCOAKtT94XrZnA5BE3tUTSKeYslqre646U8AMM2njT6RSgtyfdVDxio1mnhzkPESgudLWcK
oBfByXmTojcRzPF2FbgUp0gyTtudZjcj1Ey+R/W961miCJabppCg86Y0rkH/b6GKRVmz/voJaJd0
WE4Lil11gIWTupLzpy9vm7skQ3xCnH/D9qMIRLdEElID8h9tg0pNb3DJH3ZocRRM1llpAsmOOh0I
m5+ZEPYPQj/FKsNK+OkQmuo7gDa7GQL1j+lDtbOBg4hiAcNzsycrmhj4g+haZ+q8W4Zumnp6ZJxp
GT2dq/GbZnqDOxqjICO4L61gxVZjPE29BVYtasuqnrGN29u+A/w8Pf0sZ2ZDZoOpkcoycC8/a2kT
4VhV1/Ja9XTRCsAHnwHe2d/DM9enEpDye4fkPE3v/z1alaZRlZ4S/firRCUPaF4sYdyplX6GnDjB
hXHEIy/P1TZ+bmqn0ENnz5SwETi4d5Xh9e62Q38Joo2uKer/C8R+U9DFxVVby9jQECwfwy9i6d8B
93WtiiLkxvAD2yu2L8UwHTkyJFzb0VBAiZehuG5By7qTj6wKXVZlakyuEgW0fxEgUxdlXELojF3f
z206orzC2eXTdEXc2o41dbfW56Y+6Q0pHMlwez//btjPhUgygj2RoDv0gpGisLq8Y+nEplRKDT7c
h8cA06Sh9k1ubuJAEZJuib44fm5/C/ukSasrDGLlJUmNzmLs0kN7yUPQum2EliWqWyNurCHazNcw
nWbQWX+o0yrv0TLPsU08ncMPV3fKNh0X2m47eDDIa6/yVpN8G/UWcEW3pwfy4BKyV1bb6iDiWarm
sFDPR9BD4DBBUoWe+jvbAHP6wghpiSLiy2uYba8q4MAhygZL/DFF46YnrZ/hwAnxD2IKvCHxCeZQ
ADo1+lUIRKpYUp5RJ6CIYdzHzENpTuO92KDCpy83at6ZLEt0thB8IbANnIVEASi1AyKAc7F5KWPO
TqMO5daocQJrma6uDaYju1kiHlbVuTTc215s3TuBm5k7zK1ynYtELJ3CsVtqVNJfARH1ozWj/XJA
mpMzNftF0fNyeyoIXhxtTvSaP6M3NfklAf9LbHmwZT7KlSG3KTVPVQw77rjVzyKyOxQb+YxS5Fdr
ThEIFSqsB6O5oQ9hhP/YvwXfwfb8D4CYiakJFwsMoUm0ALh6fB/+82xaUTNVVuNGSTRbVhD13ng+
noTOhxJSzag0h39q2eOKzMxaAWK1yqZW1Vl6KHUqrCZK8UkvlwTGK5wHMLwWf7f/iZX7uevDo4oi
Zgn519YBKqBUxFtHc8ZZimfXHb9tQp0cURPGuDyJx/HJkPisv7ftGN9SiTP8cHSaPCRG9QHsSzyc
DxAra6eeW+66cnVy1Bq7cjQmccs7yQEICIolJBLBjugOw/SBLE9aoT9K038OGjhAGLlpZURmW0jt
XihOG+NIlSYmzgC8XMSiXiIh/ufhef4MvANfAYJo2P0eE0zH9RflLfzDH/3cK0OKepnYVNvbPasr
N/ZqEwPHZ/Y2i9the65JlMCPI+R3pqmQ4Fr3PFtZmxOjFCPLijPrJuyv/Ac56JZi4VaZXHHnbCqQ
KBkWwN4Mis3Xu9QMPy9DZinm9b90rjz8jIhdGWqWDjGfnKNui2N1BcdqpK8Tj6jIxQrLyXDwHibR
ZUcNT9dP6JobGOQDntLFQ9OSWwXaUEKLbDGg83uyA08Bn5q7dTPGYzCg28jaKh4WGyrMp8AIev7R
COSGegyvjvDN1jjEfJBgyAmOFDaqJGOFv5TMHkRCr0mD+o+AOyVw0sCszNLNRy5AfGHi7NdtucsU
RHln3k8uYtylHq7bD7/WZRZzfINFRyTA7cZ0enZz6xH9a7Ka5IWv3zUN4GP/5n0v/VldCtmo2YAg
jJbRQYu+5J6WGpmPFIDWByfSWIAG5jrL3fgfOrxSl4pozxLEZei0WGRTGBZqgGC6Qr6/mQ5zbJml
voEVDxhFzcPapC8vl+5yoZ+nnpuafqEBXNHhmEkJY8YUViYKtFU30HLZWqFVSyjpQooa83GPeVwH
bo1qpIbbc995581x2C8FRprJkBKBkitq+I+PEKRgsjK22b+nFHX45symsCsIciZeN+bzdvAVouHz
MnkXCmxLNyGjCuMlfuTj2xzVjXZMBtuC6R/H3uDVa9ppaQ7T22mfohFZXKpL2YYICC0NX1K+B4Vh
C+NhVAfUpeg5TjP6vTiFTupuEGdv7x2n5G3eevckYF+zrhOEESSDGtHTKFBZY0j/7em2OUCSmcHi
XoKAIRdWtOPp9C2CpiQ3kf0S6YE1TYu3pp5Wca8q6WxCKDlj0zjSpE0Z3F6dDawsJzWj5lJ2n61M
Ro2BxYCHMKcdt0s2YtlHNiYHij6ZmKyjU0D+XzAJKcG5sA0r2I1xzce7/0+ACJmdrdGnsls5s+2e
fymWVnLY4UmU9qH2eLDJoVaaQwHcx0LP2HbUKu7H9KwKD9i/tki18rK9g2r/Fwi1ONll8TisNkel
jeSuKBVHbxOLfFpaByPFrm78nTV5D4bxbZJBZhEeqDK2g0kGNk1VxlK6zXi0m97ZP+Ovq7p/uYkC
RlJwzi9ns+9mKFX+rrUoe1WoQjCIww/bqRIpUcTnabp8w/YTZjWPj4U1dIvf8rn4FK/EaAvTMR05
IMqn+ILhTQNNIkOkNwcDPuAj5+vXYMp0l9GFgTjnzFtI8s6l0TsBClQUp36Ej60JZtX8cWAEZxIg
8/EIgOtI64tmmxNuME9KRe++bpcbg3qZ6uV46DHaa2/U6CLOtfmJnt65/Dr6ETqfQnBhlC3kuRXY
qvG6vJ0jg7E66Lm8nqYal9tRTfTbavRx1hWygHOxarD/gPob+ssSCEnF255MER3AKSQdKpatCxpH
hMBRP8wPV89oYRuDpG23pLYZqxlcc/cbmcZKW/IUrEnYB0XiEkyw1Tc+YGnGbbLolS3Qri+56JUg
llKHflO8Cgx3iThZAwnUnl/M5A6/dWUR2kgYe+Yo+vEsYDSUiUGw1ICq9xYI9jqwOpS2yuQF3LFf
SUY2n8R+/fEVcthKCN8zHjNaXyHiRPx7/iQVWXKeyqG75FlsVOtrDgytKVaBNqFNRphbDM8O16AD
dpjDwP9FgMKu/FUQ/Raq0H5iIbGzo5DsiyACaiiB1mhgVl9N/JEl+gtkVADhPIomWW8jaKi5fgeC
eVyZt1fSckZMUDADMnlyej9xnTJIJ25HWGLjpMnAt/L5sBjmM40F+jiuCfdKiK3GP3KyDaMif2FU
BAAv27hoXY6dmxCyqN3r2X/blpoDSRX0yXWY8ASI6i2tARo9+MlNhnoHwYXEpzU5Ps7121hImOc/
Hgay1AoLOzV4IdCNB+hLlv6N3N+qX/e/wm+2tQ67JSr+C+NmWBCZlEuNCOkoO+X1SrTnh2wIv1So
Vm5+BAbXsfSaX2lxYKbbsnAOogNMNOLr687G6jXRQP56RasVvjF1XntH3p23q1GCbdmWEDot78C0
p8MghGwpweCSgby+niHOGzAFWAoTNJeitorfNOfqbgAKv6fsRPuY5x2RLamY/rk6Ii6Hrw3BbCuD
hS0l7cDd1una8fn4/AJgTH6GN6Ee6gz9L/3KXb13prbPAYRdyK+6Z+teBAti/Oh/gRTtNwA7uxMS
ZN+IX0NmNi1TOr6w5T8+VEZGRaRwlkDTNjowpZtNoHyZi0z2F9cRnKpSEjNa/bLxmlSjwqUIZfeh
xTOxCM4Rh9z5IHCHlpRj/Lp4Q4jpQK4H85r+LmcfqDZxRFT4nprGFTz0NuzYaF7pJ1+6Lv3o6xxl
XfjzgvJhXRBEPtiM0sI6cUOPFBxSlifozKZwS+H7G+G6Fvto2OU8m+3jkPnEZA76FinvitCwInlX
U9CADaRftHDxg43LiVjXGi8bput5LFmiIzzpGHxWjsPTTwo76D7Cj4VG39kI1NWM1IhH1Vo5XDjj
025OZEtFTwclJ1SK4mIZw7dG9K9XDlI7xfqPMxePPrHMTKgigROMdaJp893X+sftciCz5kMLsi9G
Us5UwJZO8FGIoZQMGndfgrjm3Wh+Vj4/i5CPb+lns4VTigvvMc6DW+6yGKfzjfUnt+ryLGz0ChFB
dRTh6rPAFixiA5eEYqFeRjPYuJgllRDDOB6rtfl5xSe2+xHxoo7tU2nyBoTGkUw3A9F8hfferOP7
N1Y80RqVwEEBCi8Npu446JN+YycjWLqrgYa840p2Q9sNhVf0m1A68OaUZi/U4FBHFJq7w+E0JYnP
eBa5XgDGhDHSMHhd4mb5s1NSsjeVBuypXnggA5xSIoS2DpKNFApfhoniiYJsLQYCOGuUOxd5PJdJ
QuBlK6EKZp6Qg4TN8Cq3ixKUCEYYh4mc/I7wL+wwMpEOCF6cIHPyfTKAgdD4YL7sY4C8HolBCk9C
Zi56fS+s8Ygh6o+pGDs1683lKWZdVjbup/UTQtkR/W6c/Ptfkd7FgmxTPz64RJKD4Mc/TLdopSBO
ZerUIFWntoFzueXQDyGdggB1lb+6CvHJaU4YFij5rb9e8E/VlcUYTQXBJlFNBYCG+zWyNOq5xS7o
+eBG4CPxDb8rCxGMux6Uz2uNuaI+Vx7kdsyAzXkQA+yrsWQFqL1Vo6o0nAwOgcOduunfVwE/c3RI
vFEG02xG5j44aEHtx6Z/rb8UbvsrDlcy+KYomlnoW3Xa64fTl8+a1gRuKsfNY85iccbagqkPOo64
QPUom0BMSjPxpXxKdjmS6dmwpPZ9e3OjcJZkAdAB4rqjySAmWNBabne7af7J5ZD9qvgLgZIJAgH5
Y8kZi0uzNqdaIctSKeTA67+mH3yE2b4ttQkdtMXasXM+t50Mzs4Jd28MgGUwBS19E/Rx5z41TWj+
/+F8+hXWFuqPIxv2zh9fdrt3Pd+aUi/WvvNjxgzk9iHd+rOA2+cBrVfOp8KwpzxLHhduW4GvlEMB
7zDA4GRlk5Fc+7d8k5iXfgwH4smGEyzsWRL6ZWmokLnEKJ4/QkCFAK8eN4BGvXHOmRrcfI/mzlyJ
qklmKQzLU1O3zzRtqThCMXnmaWgJuau4v3ovIdRSEDbBI3N19IdnyefKffPwSj4HatLlDqVjR8bp
D2U4ZR/oR9fQdNO7RIa2UP8AZS4tJ6l/OvaNC2vXerkIghMErBDHzvxUplQDVmlesQCmnyqRyX6P
F45MDS1lI4dohglNGDIj9VPKrTTMBd9czjPKt7Bchq2EGiHQfiSFPkQ+vMIs9boBjXg5x9XHLSRM
wh/p5XOhwycuRyJ/6kTtnikIbnKH9XhLZBfZ78CzhHUmmwmFy9GSU21JlLr96sV5NDcSqxL3oMvE
pKVNrYIDJSZairBoK0b2RIoZYawcnt1VBjRoJ3TJIHPmRGxT83Q/5pJh/ira9hEacsUECZtMnNxE
m8ddPTqVW0h+qO0GoXZcsOrN2yfWT66xk2J891GGlKfHycMtIgeqTMmdJWNTBNioUJmKvekKibVG
fvsFYFhC8f8CzTvoYThdZt/BdWQFcBtaIHx5FytlQJeDbN1IinIuE48D2DS0FzFrmnuwiPBDYp59
c873HuA00YsUogCT1xXFf52NR3/TY7TAH6n/an5bFZ2097nC4sjNrLeC57OfEFBZOqMRkiv+F9Ul
/3axfn7oTm44QdYzvaIuo/f0xLknMdVu57xUnrMKgUiePFE7WoI9ZqZhibIaV9fYbtE58anqNY6H
zIAoQTWt4IKASAFz7xw4PWYPOk1s0w7J6TJCtDGsX1LBQAgdUX4IoOyC58JtzX3DkQ2S3YKyDbMZ
1Ip7aEx+RVYcdHGvcWl5yA+Z2fNHXs79pPkg4fOGS5tsQPMOPidKuFXlOHI1ldzoBL9+SgRzAa4D
qejtxGFs3W/5OG9r5AMYnuzfSEN42GSAR+FtM863CxTxbeXQu5Qtw85T1WK+7ydWSw1ucTCPmTZy
HHQTF+ItrdAfYSiXYqmfn78+xQYk8kp2vz1KcwRQuh6ZNlZKaj8Uw8uGkg/PiwayOwaDVDCgKsBD
r/Xc9BwBKw1qN5XA33IjTfelI78CzOurfkF6ShfsbNLSulC8L7jl187cIxoUNfKkPVHgyee4Vm5U
TQjVOXToXicLXYedR6OGVTdWbA6LqrRq36TjJhEVoEODo6gSutATkFemEsK7C7ZCe7VFJOtsSYer
PynS0LeMMBYkyn7PkOYsh3WUs2Dx5u9LBa9Dq2q7yQXfV4sWUXpsHSlpqGTDKfOUNzRtmPzUAn3R
nbF5HDAwrtAd9FJ6Vw9tK1pDmRqqnmYT223SM0SuLuVqeSQNn22pGwLi7T5ant20117vlIxL9k/J
B23W7bV6euOWbSmWBFv6Z/1t+fDgcpfjJuyJbfCb7y1bAvCJtpqhuT0M0iDFnQdyraS4YbIdaiNA
JYphWcr9oRUBR69aYbAsdWdH8TQoX2VTwe9vj/eNidUebeaWi0uLHFdpUx6CK58nrcZfMghQhYPx
0KaeSLA5d2qiqOAYaWAgIixBKqkFms68GP6eqTKfw/Q7J0OzVWuTZUYSHkp4Q98hFkr8QNpLN+Iq
3UzNEqloE9ME40Gzo2ZlagcxKU0U3gSPHNp04Hl+Q/3kgVuFXeAXZedwZ9VcMGM6+o5oUkGu5T/2
tO7mlFXroKy7to3t6kr44jNBlj6IPcT+jeQYe6yadligfezuSOtamw4bwfYWar+MjPlAExJrRojj
Rv6AnVC8z9ybjlVp5s0+W9EsLjwVligbkoe+jWn4n4D1t+eTjEOLVdYOETF1V2sYqrfZ1NAezo2a
FnffMsRTsmz/wW6Oxt1VSvILQG9ElvbCKT1Mb0qFqR9myiFKyUzz/ntiRw0K2CuLUc/j8Lfuyg+M
c5j3e9pCmbIePnJ6kra+mIw7sWqosG5fWoQfkh9f37FBa+GXDmkZF3RPZMi+GAI/FI6y/U2DAPdR
kzhEXFeLw4/TFPogprvqGw/oJAYr1COjlQjLxbdierMgAL/SUOV//BogHe0vUXGZVAxilshbXjt5
3IIHjyTQ3V/K7VvIyg+grWIBfxVwBcy2QnCXLidwuZrViqfr2CjMkwwrYhzZA1kmPLq31nWfBJ+O
RlTR31yXlE5Jf/Y2yqgdyHoD9TOnxcIQB4OcefGBxG2hwVZVdrWzVwPO0WDKLhk8OMdrH7oGfwOO
rMIApoaw0+jZAV0UBPGxMwO0oh3Z5rC7DPmzrH80OWga+sj1YV3TmkI2g88kiYIFPBvZQmB8WsWX
/Ka4gcFr4r0kRWkn5E8mk/zavc1WMiyoojgI5a8kL2ZmK8UOTpB9PtG+QgBIImNcnLOWpbpyD76F
F8I7UYOQO0CdZgJM9ktLR8oq2VCLRW7OzMlTj9TETj0Z3EsARiEDxD2RbrlfI1F4ZLc0MKBJvA4z
at0dCH8mR+F+xQ0MXhOFFvwey/8o+KhdRlvkabRM3W4mab9VvP1lHo8LhDvdXBnEBZyl9j4KR0b/
/2L+QPQTY2tJABPsSg6yQFv7Y3FpWgBuQTcScSv+onlFsskme+MXMsWwpAozdGkIe8WRwMfQV+Kw
Q8u1+dzXpfdGc0attlUnL7rYgGDSH+g0plhBNzMkQanFgmyOg90H7guCY4msUs43jLPoGdCQZUOR
mQiQohqqHebK7wecHCt56wkjH8oM09SAukHg2ZCwtdl8USm4z/e0E9GxloVAnMYijfTnlfoilQn5
BQdd9xnaVtWNKUnBJ1USQAZz3MD/3tH+2Dxrd4FUPwgrRBrHjAi1eNw0LjPdiFta4AwngW8QpkwB
g1BumdJSEUoUnrvjsCsoRug3BwpgsIVUV3lBAp96MRYiXAGXsfJOBW8fy+qDrShqK/8Eovw+0FBj
AYBt3SrU5T/yR1RHdTmoPXp7lTjRO5/elqSK0DsgFo/zXAX5lyT1mfrj7UfMLEeXSQ/jQbW9mDR6
pfqwBShBEggQtI2A8CeKAru24k504Li/rW1hIJ5ZdPsZknxNm02qTkSyf+oxpNQEV1T5wCe0ArM8
ob1LieD2R+KQkw9TbTyjUxasylNoU3Y8cc4U0hGv1hPRPbrBkDHiKOT0qgequkcsJybeWGH46qu6
JQg0PveZX2zbdJzX1V6PC4N2eq0VOdnY+DmxD5z3OBSzSq2v1YaJ3WWg3A5uPSKfZuLrj38rVP8b
sWEA37NuhLSAjG4a2fd+UiWGF3opolwkP2wHB07U+yaRa2ZGd7/BSjoi+ERy1t0w4EY/QYAvnOQB
MaC8YKiGYiVzmNgC+FCjJRYHgdH8iHGykSqBaO82sAtIMnwoie07F1ZLJyB7lkLrC5szKHprBhgA
st5iBVBGLCTn2IP6Zdj+UPmcZ6N00I/yjKTcAkYEmImsUcYbkk9tLkZUdemUHC4uH3YS7VZSNw+2
ypwbBMHWAMfXNRd/IVVAuwpqBPASPteuxtboVhKMUsCBNCJ8PQH05zmJaMlO96iv5Wv1vX+NnfuS
eW6XYSEm4B15cxLi733WfA37bdwzBSHaseaDJoEUATCiY1/hH8GEv0SuLWOX+4qyAxEMaI6foYDV
Nv+T1DQtOIoSD/7AlTEiqU2JqQD7god5UeBAPFBhMXvEhMEnXWhihyLZJQw0l3rjadSCjlltmAsp
TGTw7jyq5zcwCuzMi1eJwzCOZLRYqi6V6iIu1IJIm9+/lkts8EJtE8jB93HZ4CBCuQolsbdbvgY/
uZl+J1O5ZBeX5xhfm1oaO0J31bmOJGowjUeKkFggaKMiBnijLEbxQngp5X5gZveYFcvPGfmQBFiD
7blbXgi027mL3cFH71MABUguyMiBJCVKM7cWrqUlXL9myUfBFPXiVWvJvlir0Zl74U4xFS3RxO+w
XkLPpNdD7YEo4Ysly2UmDt3S3VNZQAcu3rpbFl0RmPYkDWVNZgNbFFDIpECNGJhoLwiX4oq7YmGx
Klof4JxIu84zq7uZN1GmiMs57pZgaadMwEX9WgwLV2D5C5Y47y9ch+1ZC2mPvO7jLzUTocUse2eB
MF0Q+eJ+xC6Kuizv2X9jA1EHYC1R1s7c5FJx13GQrrQs9D4L4R52DNsbjyM5lR9pr1nLmL3tvDRC
BxWxGdsw900nvSY+3cTDlyM5Ntp9DaJ9ImZ3VF1OH55/a6QeWIq2o/gYvqfqMqeY/7ZL5HBtB1NV
OSAvnE/GMQ0GuFXFbXcBoaJkN2vIUADVyC3AeFTe9mDlygiq7J1HgBH9hbZ69kHuHy2QlDNPY/uF
uN9wF6MDTnxjkE2oYTYdtuVIGivB6ZM2RON8iPUxD81UVU/vlQyQbP6Ig9eg6jt5XjUN5cu6msAs
5q+dQlUgb1SX1gF6BIQA0jXl8GNPfSq0Xy3I1LMgRSL7ipnLuTvRrTtacuAA6yqH1jT7JZHCtdsO
G6ucvwPra/Szkr98cK2/TPR2pvePoJnaruOjAHa0JuhdvC4sxm6s/U5sY4nYVHBkw2riDJkRH8tG
i4GYP5hLX+dcQa9B0tepeLROwo0ecoSc0kA6tG6xbuQi3UX51wXpkwgeu0bym8olghQsVpKcKuZT
B0iSyyhIvzjjqyRwTcCxvPk9jUnWyuKgh5hpHqO3kIzBj3NFHO5MS0RF6tkY6v+oCgjq0seHswsB
7PIz1P8S5RuhuCJUb8GEP27Wl+DzDFFS01RBmk+L9g3GXya64GmNMupvyxjOEjgo6WHY7OOQE26b
3P+u3Vs39JvAAN5kZwme7Wy5kYC78nVEvjqxYRe7gTI0QA6GEDGspQ4io0Lw2+G6Ub2HxOr6pIML
p3KZH/QYhrlZt0xI58VGkt0tfoqi5RDBA1Znmv1bQqSw3Hf8ol0Eu9K4y8amSvZq6R6bruILPzk2
exKaHeHgddmyPv/IBGD0ectUAMMEYEy25afOXym9xCzpQPXjCIU5H2jtY7HwzdVSLrpg7m8u9Byt
H6TqOAiL8gtzRpFbUfzaKySon93aLaIY4wBIhEToWgFWIGaTXJrw9CkOXN6aP5UE+Ymxe2wY9YRi
SlWIHeuCkeQ59d/TrrSk34Z7Cx1uMRMkG6vZf2Hf93EmrwKSJUuw0KlJWMnkvUS+tJKjrQk9TS+U
y8RROjHnl2f8eLZWy8sE/D7wz243qGmo8VorBN7we4uKzvkxdhzds0/2SBI7eOZoIGVC05eo31u3
FGrrvKTTgVFbfz4mU/otURK4rMm3+S3ctFzjy83OMr50vNQXjTtZ9/buPCYu2yqTAw5aMPi9V090
6KPyHWOQCzn2FsyQrlaHUPLwffG6d0onE9kacwLBRoub+JX1jOTBJcMuO0tDNrJsF1FNPKhJeqqB
00h+47BIFXQXTmjXEZ/V0tCNwapSzWYmBF+pj+N8spWgzzhzAVkU3YVs+WqPm+uNU95HM9OU5Xcv
ENzq1bhQg2JgJcePjOulgtCa76qY2a87/m/eCfDnxTzPbUPIMSBDswEwjsy00YCsgfpJR4K9BccR
5cG3cOn4YMJvthjcpzwaLkQKA4KW/sb38GNRey+CgXhB2p2bQevNjNKEcVhIVjThhI5jPJqcaPlj
fiThD49RmdR/j/jkolqPljp1YG+JrbKpclPCfs2lxLq4+4FyBwPm+E0v4k7tbFdN0MFqimhODYjU
Nqup5ykZf/q99+Oivgoul2jBL6zKkPijnzyDV/QWeDO1CsccnYE0zCdF67LfedMb/gvvJGox/bPC
zHyboaMXoEEQyQ0BM9QztbloZkiUNSFeku9v5ijTVizNY8NbcIXFfmfeb+XSLZtbtI1nCK8AdYxK
PsuU/0XHe8OGmPUdBmiCjWjEjIjmIAOWkCy08Uw2Ga+0ao+loVuro26tgN09LwX2owapilHuHbt9
fj774aM4pVDbFYFS3k8bi/yIRvIp5QdKsniGi7kGDD/Mj+iYfmiIxcijIS6WdPTmt3Hhg4JMPG7E
n0VLjYLRFnFHnbgJ+uAIruu3d19rfoWEdDknjLiHlrqt6v981ybtL6OR9inq/ymzrFZwEaqcSUvj
/M/16LjHghhSspIIntDXbDhABwFcwwI2lTFhRa1qstFpb9ND1VtmQaFst7t9NP6yXx7gRxaV6szQ
gG44A0hWmKUiLGJFbzcrErPSP403PTHEMoVVeWB5FkVdrQszegMOOdYAFMY8rsMclssi92p26bF5
BSSwrbD6P2zpHd0P9gauSE47eCQD8z+SaU49MykT71ZPZJUjbFpsynAdksiTOMYXONOfEsWMk8Xs
zkHqYxCqWu2sRPg3wVbeA6ZPa/8DnDMWJfmjR/xqjLReAGARYqL+HY3gVR0z6VFTrhwdT150gFn8
0eWiqj4geiDQsoNRQyEl5YvWs6oQYddBK71L5nZK5ZsquQP3ePSHZyuWGraIQ2aZEvmhXZbqJ53N
Er98cm71J2GjeVZlhZLxqiWb4SapzjkTOfQQOxUOaiyqc5l2lCdY1BxlEED61rh2bt8zrcJl1XcC
vrOpb+u/M7wHRrdq8isOsUwxPYna8+YPeSLNMxPJbU0AnUxpaArOyTK1/tI/wLREDi7CM3NdADWp
p8j9V7gQxuic5WZCfhFJ5kDp1fMJUOrpnNOZCzxJpQ3ffTLIVN28eiVM/+2HEyOSe3BJhaG0aWR2
GMANxBGZXpcusdPJXeMkUpbFBSGbTD5SaLREcCz2Emwl5Nf7pFf7t/2MzV/6+eoWlgNtmC3H2ooh
6RT5CG8vGECf8DsgZrdgWHvX7esSroEEROp3Lt5wXjf7PRroZzEajH872TEtCnh5Im4G0PZ/YZqq
Inn3vaEwAHqBebDLWwpnMrp+lqZ03Ilz6A0KBSVEWezFwCGn8Lit4plapgll9S3AjbNs4R0vMtcz
U00m/5tPalMKeCn+R2H0i7f2krVe2tGNEClQ4HIYzLVWQ9iUnNJA9QjzPtFsvWW8UguS2BBHxSa8
8+k+qn5nKXAnGOw3GejlOqF+Qmbmpg2mvj/TndPDSiUF412gJSNROgySXSzADITRqMb/KEx+LCvn
dvzYgLtvieMiSQ61CBlC3rub+FrDN0xq6HY9BPJ3nieAeuac4+94wO8l0W2Nh/RtJwk2k56qKdtj
WW8fVwU0E2ZpvCkkSttO/KC7Hake4QVyeNH0/PoyTB+b1rBapyZOzSL5JgmLogYUygbhNR7qs7gE
/ACqtKvRDsDus/iQyFDP36W/I8DbAz+cdS4LNIR4ol9bcqyB/c/TcfQ6304MesWLlt8oFoIbYN2s
1f8kgPJpwFQY+9GVG7ssAJGe2yE/o05xfwJLnHFtxVbmbR0RF4dAHXRMDMR0i4mTSG6ZyYyck5pi
OXGr/xOotFZZsqgv7gu62K6h7uJ8ZVTJS6Dgyqe3AvUCTxrVCB0PZp+5veCwknV2pyjQa8C01EGs
6X7hLIXK3TJ3Q15ahLx6Uiaf9nFv2hqSEH8ZBSkkK/dfElvUFx8obluXmjvFC3DlIQuNJ8V6tuW4
WOyhwUV8Siwn3fOnvxASYO+YO3u/zqcEBUwH/UmFJrVhdvI/ZKpzhJCLbaYUDK+xuHrrPuYCA9yW
iaIxJFvWj1N9ErwSBBa014uws8Y/KAbXV/egDqoseCZVhwMPKA5ukE/nzQu3en76f8ORivU05bR8
p9Z5iUFX5GqfDY1/39729/ZIYQfKDk6Qle6q77WTVnUd/11HIPy/WgyhsWxUuc5f+Tkx1d/WC8dL
B+kuucJrM6zwm3tuiebd2ZqotdPs6H19WQ3zda9HGUuwZhtmV0ztLno1eDniL2osFYVt+tEEYbtx
GAVMufiVZz4Tuxnj4OPjYC7z7BB+0svuUwoSd2jUF9Pms73qwpqylnjOm1r1ntJnpkqpPVl8jvje
jP6kQWmZANMNzOWsSp8xJYGT/wtCln5MjRF5auei5Bdg+8QSMEizPr1m9HkSVbgM9QqMhiDptEpB
jq5RZvisk8I88oCcdwo0TlqeLbgtBFPHigWtrtOpjh6eLIHAmhzgTunH2HOTklUXYeyCtad5pyBL
ycCmp0mwtEkSO1LpjJcL6D2DqGZkk0H6lKzFRa66SyLl/ZiQONlJ+rsrp3MRqs7EiGBfty8X4x47
svAo5NEGm2/kXnTIpu1uMoIm/In7vCoc0eK7F8Nz9rb3ilR2wt5Ybo+pTF/F/3IvHULYVxHUsFT2
iSPwssOYxHufvrW1dO7fIy6ZzWA0NmQgCclLmnaKM2sdDerOmO1zO0gJ2XHhE6dPyD5UAKWWWt3R
MXv/qR5T01EadJqfEDAd6X/q4RbqYPgz/XYep6dlbY9TMyfm4EWa3io3SLYHyoGJhKGBYSXwuwMC
X6318yY2K4gS44Kk7T6C3xyR37loDNO0bIYJZlVnIM2jyS8hIWMPLgdvVWneaZINqHELp2LhINP2
UssNk8vs+lx5NqCpJUcLcz3RUqG8bRFN9gercTb5LKJxB7qfgxrNdkBQ10TAuFaGGlcWYqvGRkNd
Up43d8s+Yp5wyzscV/b3C2weAYVXeQwZvx/yORS26qQyK57XPEOKiwkcwtITDWrcRwz+NiaMl7BB
8dTbXQ6x62nj343GcYuEt7NBXPPJwmDPTvIR7WDzW4GnwCTz26orLBikYsm5wLaLcCQaM9AJy0qP
BH2ct4LZpKEEsDxYJDqAgUtX0hms9kZkvHcnQTH4f5WnYxm/TsCO/c1m4h28bmKd4SUj5XIFN2IS
hnc14nyWoyQWI/+QVhHtbyQiZcJEmb3SLmnc/6zSx78V3K7gFG1Tajjl2U9Jqh5FJQyYW4mkrvYL
DImlLtO8Gn7DApW4eoozJLizrVVgw+vzFCRlrDbbRYhMMuJCXrBW/QGD2K7aw5jk6u06NrPTEO0+
KMKIBJriaVSw7EI9kjL9VusLPOt1pVop7ZnYqhjiHW0ZJZePUjqdvqEJemh1/11Ix+OdlLPy3Kit
4t7oypHaShNTRq+HXvBtwpE/W3j+QRWyCfLgV6+rkxgUO8roLj2ytNwaNKJFuZ22z6MjZQeG+yEA
k9jfcJ6/j1ClSzM/yz3SD6oWrsqN2Bejpnq9kys+CLqF+4/r2EgMtjpN9Mbz6f1oR2nPE8C7Dfdn
luRh3BifIR79XNohkc9IMuw+PXgjZ8YYJYXniZ5XbSIH2RYr7gsAXXIBvEv5dj1kowRt5XH0G1s4
usqQmTOJ81Wj38Op/eYm9WuFimKVV7eyUOomt6k1kVfxePXSJhhX08DCSQDnsSEr6Y70i0MKNq5m
usq/c6lFNlP82uzEPrn4hnOU5Pfd18sj/hdjLZdtpZKorGS/1au53GZlZJ+ztqoV8v01fQ1v2oTD
ZkE77LgtxVEsLK31d/y7MJdqfu5E6A7wLzns+7DOeIf3PZln+dp0NhOpPU5QlHi/ewIzVsWJU/d5
vYCZhA881sMCKb+uRr6xlehObiJWsmW2xqKr4NfitNcAWQMabUvgkk5QET3psiWajcXrimU2KsRZ
o7PhpFA8lSQOx4oj4MVAe5krbaTINM8C0l+BUyaczmO0vvXtrVHa8ArafkW1pJMVlOIcMp3/ymkw
VjcknQL/MH+yY7ofOUIaGaL6NWYWQ1kABAjDNM6kKDs5vlCaYg/bmgk6MLRcX+ZN0PhItO2wit9S
RvDVcKmrPqCLWvXEa0nf0MmKSrnzcrrk2qnO+qDdwe3NN+VLPbSOVOB1rCAf/OQdlrQutRF2ZctH
pHshtPeXRxOmLt/2U75WQAkY+eRzM+WaY6tqoR150qCurrE/D0WLEZtH0DyQVpsMRzSWjHWuTA/b
tsrhqAxAoRnBiy1CgPZYGwXj5hYcyjrvmZwDwSKyNBmjxGeYmOk9d7M6kp3/YIL8wXzWkxGGmhnf
QeTYRsdYtC0I8YXCOuyBdA/mEXbqHkFUECRYy5QNO3dqSltqFSwIoql/HH/xK6T8Z9eYHQeCA53O
8nSocYbDCYN55VbjFp7RmIDmRXRNYonTN11mUmRF84FVneHkgKPqgXHfzED2xSsYJ3zwJ+VJ9pxv
+OqwVsRgfyH8Uy5vlFxhZIalJ1A4YnuwDWEu18TrE/iqm3BDViT6B4zj0OfoIpQMojLT9VSNPTqa
OMpsMmmWFD95Hdh0wtkvDhzhpuqxGgdLu091n+7Mjf0xbYrsIbJWD4kSvgQgfeetwLbHuJwZo3WM
Hgax+dW5C7cf0/0DP0B90jsovu6lbCX/cA1d1sDo3teC0j+PbRn4Wl+c5Az52n4Vwi29PBcxcFyY
oedJVqapmjfAj0Mla47dwc3YQOl13t++XPuH87VZA52ZCCJqoFFZAa/BMsarjbQM5EPT5+VNYqcq
kwVQlxzsvKNCdbViInCffE4+E6HCNxF/KJ10yNCghKOhkEFol3MLZgTWxIAjN8DU1Eo4vOS8nau4
8nE465H1dBBOx/9PkQaqYdTyjVaABi1dKelszMxphOTARwQu6jSvjfdTX+OtCkSWJQVWNBmnG3CW
3nokOzObia81Hg9o0hGZgYstpxCHTEvdkR1YdUbABj4rCyNqZO5VMl9BuB2UkKaVVs2uLE4ddQVn
P6TA4pdJrRMA5pTYQiJ/AzoI3h6GZ9HtYmHhHOP+J3GRtlLRaj9Ta1aMxYa9+0rzzJtCVhT71SjW
eOoYguNgXwtHb6Br3Pv5M4AfNs122D/sroRxz+bKPguMC1lZzoQiyUdS6HkRF76HywM7+ub8Kn1l
E5j9qbSoff8/pSHH+WEKpsbUW7EXFFFaRalIMM4H68cBn/WDjEY9sCQQoBztrsf+v+3WhmEGglJ3
pEPfb/Iach2fkeKW6Ptwy+4TCqIJkRzwtiHvBw/vbvp/YF2cfP1iJjvtJBxBQHWTgAYKVj8E62Qm
RY4KSYK6rp+qG8S99AjU7MVhQBzTY+0ABi+QIPzcScMvaXnxuS1qREdgGptxzXIzPlDeRkmLLAdf
7vOX+hbh14qVQAwxW4GE1VQKlUfvcPFErXAiATHjNPP+okMR6XdMgfeimZay8tJd57YJW3ExkY+G
yEIi4P487/fypSbzt4+Aj3UvkLqT6Z65Xw0DhxcO88flZDzxfPuyeiVptCkNXJTXRkXBhioIh50K
IjYyNuUeO8pG577sAURGDCho+BCa1tqIWercw5mS67FM+a1FWhw9aFhZkx5eTAu6EstZSFKyKSXR
DpXefum9zg/Ztpa32Egscz/JWv1WrnhpXbXWXmgwtJVjmBv2gZVbKFJQfow8hhHI+6RhZYQwZ84t
l86O0sqJ1qMcks2LEJrUkGBSXROyPnUop0PN7INHxQ97QwR8EiWOldFuyz6OEZXuXQLBYqNtUx3F
77HzE7eYS3jiAXAqX6QPVe/ZTGSQsldTxclKJU9vI8/Q4yZQ3g/eWn/qXeKaiqfoZWXjFj6eMO0j
/nFKLdtKfbAoDjcNyNlKijcIHQ0To4olC+8vvSPeuSbaeCL7D/7B6+AnJrVltr4Q+cwMHNC2Diw7
DY9tXGKGheVw4L8K7b0VcJys9YHJGjisoZ734kG3uL+L7P+qcMZKfdKLGq7Zi/fFGlILXa4AJeuo
aoDGZAiu4QvimnQVVw/ANDenKuv12oaAVyxvpssmk+IvN7Mk/I68wriAWRCuu7OmDCBoHmPDTumT
JOh4NYZwpfNIjzs2E09Q1xZth5Y0Ml0VlMX52yxZfT1rGrUTGc/zPSKgSvt+h429ar7YiStMIlTV
tBX/cxP72AID12vvVE9tqz/lixnzAPQXnH8UN6kwgH9OESNNyUg5MadFAhJpZMXl5GS7LprN3D3L
43mov6KC3vFMjkiNCCodlZnx+optkJDx+Adi1TA92UWxS9ttinlkn15owc5vkevLRmDV9xUmbHh9
SO1oP6UPiO/oL9N6n5CRCWva6v96NZb8X6MeoZkpPgwMZujQW0i00J0BmWyIx6Fqu4WYqVcuCZWK
HOJ7JaNs8o+psZLiuYyXwZpgVJJQxafJPtPlI11GT2RcAY62ks3948Dg4gROXx5yPJgZpTQPc0/S
CUXfJFU14aAV+P/nCn/emzom7AHbmiKDUxpwv9r9+Gu2ws/1t2BpjZ8nIppYjR9taWbpbHcLmewr
5iGoX+7wpTo1rTOkpdkyZHSYZ6vXXHHsrCA2Lq0WEj7YGJdKJn+tZOVsu9Q7rejxdyQQeQ0NH63q
0ZcBH0lb80+ci9zytUf9m+m4kHd7MjOOgY7H3W7rjiK2UV0fDfhv/j68FrW5J7J2OZH3rOaNoane
rKyhu+0xZwdkCuY9Kq7XtfzoNcoq7W9HwEZxkMI1/1DI413v3dFoNxCQZrWgE+ovdMq7T3KcadQC
lH1Qg+qIqQIYpsXWdMp82aJLFSa1PXts52mVisFBYUGjUYx7pg4YWLHm+VEGI4CzNrmuLGXSV4DQ
trmqaAMwbmcidCf9zo/m4kwIWHIDOUZz6GbJtLUlYiDGVGVUmGloiSv/hxxEqfgsUF5gvDY4e+Kt
+iG9kdJKJkbRYBP4rAs+6DFbnytydr/rYPA8YVKuIY/NRSPOqIo7ycFg8fgKNmsfwPBvd/2u7eUW
h2tLr1Wc7GqLzif0WqNBHMk+FmvpGUGskLwaZxd0UWPnKEYhIWYIPffqYudKSVMjeIz7o5BG+pgy
L2FabxBGs9OHvRsF0UMzDbvXTHCGHlHy/81o/Ro4EtNPZQiG/CRGmyK526XZEwS1/J0wOfm040y3
Czff3l1rfffMqDNjoot6e1+nosuT6r7nfCONPkOecfmtTP4OrtOA4aYSde54+5nHV7nzsgRxznDu
unF9j5Li6fzhqxjLmJbfJethF9BltHcZdBwTw6vOKAIBA/td9P6xGvcIGAnj0wPGdfUmbH3z2B0t
eJyJwZycpY0wZPw4V5IQqD8y5to0bDtD0luajfF66Ioc3L/wGg7WeN50xH6+mC8ugi0ZUPDR/lE/
GZ8I2L6zB8LVrgrwaaij/i3Qhuy2JoyZg81w2PlBXTG4R+VyJyNn8UjIEJnGZvU7mlUZV9bl0J/g
dx9eCTSaYsNB1Viw0j3q9Nbcp264EC/64klUMWhORaPW6tscfBTHjtNsK8i7U/WeAqChLcQCJi70
XMyhDkgUyxBqR5tCMaWrnVO9JfRw7bLYFYaFEeLT4RQHUCuRUfcp0/JTXxzPBjXSoKep6HPmk0ig
Xzn20QOKtFNiIaXLbyOxt57Vrf7ih3UPuueVAzPkeG2nOobPaD/IMdbJysImytjlNynuNMwjrPsy
+UGOBuWS/boQkly0QmZj6Khdcdv8888I/CjL4KjreYRKhEMaP39AvuBukEvbbRbywqMDc74FUh/N
AQypm27a7ZJ7SMD/uopo639AcxCdhSrk1hm8O9YHkpzvKv14solOmaDPHndkH/iD7dZZDRmjLzZx
TtNTtplq066Q0+JylQ0oq9MGEK6mWa9spM9/VEPza7pYo/ogKEUknDP9BIab4/Z/S2q1U6mSjz8S
8F5rV6Ckpn6oYVm+euKg0yqwoD5DRCmxjGIgrMHrEVYjsYz7th29RZrosInK8QurmIulCh0LNPX+
grRNvratU3IDur2yiKGsuYPkwp0jvJKxQQjfU5TzYrvZ1s1ql1DzmHxyC8DUfp9PakqTd2OEir8t
NSu0JIqMUh9vHA5CCdVaNDsf4lubVEtVvbtnBENgbhAMxWVmSY+ERRA2z6X9YUU1qWsWEgPBOsxE
e9byp3iJiItNwsmXtR9qE611wMmiclVE7kMfqSm0aUbFqgTTg0Tz+W3Ldq51DkSIi+7zU7Pk6QPs
Br+bskgqefwsB2FX8vWMx3DLtcD3WjdHWyMPnZ6INWm0zil5icKMJMBjOHELqd/1pYmWhH0UlD4U
t86UJWM7bV1ZQAMKSKbgOR6PNkjm16hzw/ebKm5lERwPg1E93ldBXw1H1nbfhiOXe23BEt5HPL5o
dGWEgWnCoMnDqDso+uI340+nxRW0ufY+4jWO0Iyhb4E7bZK1sTJDxokhv4fmemYe242a2k8wuIbK
f9S/ptKUELR72HBSxdSMfHhIzZxECvBj26zf2MBDMNdEamnUF14YfAbr2cwFexGMoJgPnQK3Nfaw
xssAUkFBH6lZ5Qmt8FO3SEbzacpcecEUfNPtKqYvZLWH0jVLpPTof/5cAOfbOF5afV+MNAZi8Wl9
G0apr7GAcbdzQ/OermXYuOFaEu+URG1UW4tCgsKgfB3QJJzHDShm5Xn86qfgsCWwX3tawCMB37P4
r+7zzC72vKkzFRcHQeqiXYtsG9Lt69gwMPftrSj+9jkqCbxcRMwSgSW5qE/JfNWgT8oxf61Ckbji
U4lV9pxlfPLQaznl8AzJ9wSWUc4h9/nI+9+mKeB8yuZqLP1N8GF5L8nFeJZUxo2I21FsfyQr/gea
M9xNaxi4uEv6Nae/7Bbsve97driYYQnJ3z01udWXmN0z7fxdKV8+XHAoHX+fHe6wQNapxyO/NeNW
QCdK/oTcDc7mzFaZM5AieULTP0qz3THu1TL7quDMvvN18/9t8xcgkZXSFI36xylPNPldmZSafp6M
d022xC9RTufnRNmeZfbEFCvm7q7xv2CnMDIdmNi0xlBUhSakN3poAa2t4kGweBN9FzgrCRzoIixM
tL+5slt4ogWDdVPfRUUwoOI2EHgZZKM9879PzTergYt6rUjTVvMiHZkyPnWzyh6UcVlGaXn1F8MI
NO/LSNCF+c2jM0QRzjGEg0iN12QkFbDtBPc3M2+qj9Q7pWVxKt1KLZfnbnKMqc4lo0S+Thb5idhK
ms4nhOlZjqqqJ0zpBoK3bt85xsIuN829mlQN1+BnsvczieJ01D7vuZGjCreHyG6DPCfGA5+OZwAF
oy/a9iZj7ckMvoqJWYuI9YxnrJL4UUpuq5gHm6o8mIrGPsjQjFINfCoXigm7mTRf+M0m31bh1vWI
GFBY6BOxrWoVpZ/sWBhxV1r0CIODT8nMHZxYBWNu3r1saQoAiImm3JvJCzEInxmf6ShmW1REb2hI
68q61wOASBCszX2owNdRiGD8Kqj3P71x5jErwKUUDEqPl8EoMzttrKkT10IosxnpWG8aJGWmavpI
mlxVvhqGuKE7+xOQvDgQ1Rw5U5WS/YpGgqq0b3PjbVJ0NGBpEnPe2YnDGXftpbsDaQSANEBos2hx
Ug4lDroAF/DLDIIJ6R/U4lLuqnhENJ+KNOFVNzwjWNtMCzNUf+WUd3nqI1e+oY1uadI8x9TiG6Ur
1aKfJpssaoxCGko7vdtyDETe791eOqRxZUn/Cin9yluK2aSV3NfQ+dKjyGlpebkS4ejO4+AMbnoa
1nSTKJMlhDoLIwpZOy32in03vw4lTpPa9Tqiq/XkJG1qIpVs/t0Fg9LuwYYHRQkxYmru5EUaxlad
R4r3p5RYYyjCAsG7FHvEgQnC0A3xWl4kG3YnU0z8OL4zPbIaUrUk3ueNNzb/TGeK3mrWeQTRCZ1q
NWtYHYJn4AkRKZhQpmt4EwX2hIJooPr/BFfuPz3tM5U6VNeJiQG15W/+jBul3gjDGGreFR5x5mtm
XJzVBiX3Av1FOkbmWObo+cppBUdjSfJbO8RhNKqHXqU7O//ZxcDfj41x4M2MyB9PMIUVGI4E+Uxy
aq8UbSfzzv+nG7OHn397x5Y2NYYXRYNQsfKVrbmEEUCZnx2yfjAbmO58GQPlkBKBVOcBcWQQ17FK
tWXObvC/kXc3OQZ9GqnH1JSkuSh5sKIKPdxGavVN+vREaLm2CIvmW2HiexTRumIc1zuk3uhGRV/u
5daLcysS8tQq47tKMYYIodpaGKZoI+C1xvGuB9aVRUYNJJCzS5a4D6vMnl07DEO8bBUTnzzgpTWp
1pjPlgOtPQw2fcD8ZN6EiIkAmYZz2Liufin8PYNKMIroH17vL7aB89k6uHi89XyCoeShYcpmQbZb
2+7ApsYcriA7HAc7VE8JTfs6GmdGpLqG0Wz56qpqtW3Oy8n1fsGEhMxI16kNS+/648m1Ji1+d2h6
njmb/AO3HMZzE2iUxqZqwYkas40QrjOxOFGbxevQ/Yi2PWlnLUTbn4iYXee4F0nkAyWwL54QoPBO
0T53Cej1/y/zAjc3xwKIDevBAH0kxsCtv0NIx9USvV0L8/KPPYUoFSqp/qieCDPGng8OCJweCsoW
49xGXV5s6HUclT+OaTb+dbolYyVu71ssXC9okeWmASI+NhjjS2L/lKukMw6LiFsDBRXK0gyKIfok
hB4u24S7OctHQ0v4J20LLaVrbyC4SPTCl6ZqDo36etgMZsXCJqjENn0+xgPUvzyY2/0YEd+6ZwYU
2JkeRtnFaqxGGsn2oQbnX4CfSfO7KO4Hzss4C9wO3HFIrHuK6zT4GMtqgTH7tVbO9AI21U/Xqohn
WMsyMz7w7sHiT9jiU+h/ymqNme+DDgPK8+wDB27ATE4tmzZXL/8Tkq33gKrnEKoGxHa2td3GtRsM
1Kcq46+HxqaF8O23wg9kMg3usgR3zNVolIgcHIp7NilZHFG+xgIShM3MgpqMUvcb3NcTqEiwJsdr
wwBptmXdK+aqcr2oVE1jVNylmNLFiFfQ4R0isn4igoQubE5NPUxaOb2+1AEfAnexKcgzPEJNLEIs
Qg96w9NBkRqOvPkhBHo1Jku/tSxBcU4JoM4jdV5tkU3nJGgQz+fwCw7jGciJanq1bjw2qExRX+ZO
DA7rG7utiAhTM4Hx0Q+sZGfVZ0LuCKEUr2staOn9AHS2L10g+xQLLEVfqHuPhe4+AxduzP/7PpsE
ROFPU+BYMmgySHdh0IkEalwtht27QbT410hdby+kA7VkyRxJci8Dk8wgYLisPmsIcEBSsludzMb+
ffy9WqTWUBOddZrF3znqAy7bSh+w4DQFKj/gOszHacWdrIZ+DprMItDxE+3jkpfZid7eP6cn2AVK
pfg5AtMXrTfvtJoOuLGHMBXqKJ2k9p7c3snpIpnO75EJf1c27idzuctPpppxX1VG4kgUVHEXIT8o
XBlg5C5ImlQ3lA3H2GJItvVWuVdL/r7ubRQHdP+bSwF0ELrk7lDgLir7FTXpLXUeJ9eZbl/trc1m
sGqUmgFXsc9fYJD4+OciA4FJg+abmrxFoOxbIW7RXmyQBCkTqzKrmy571I6WgmWfSjZBTPSAJenO
3P7HS9CGXAFAtVgXACNCbXaSsBcB1Hs1VsyDpfJgeBwhily7a1FqVNK13Y5x+TllbGARVrSoIbrp
HnJbmiz1vTWLX+N876HI1t3VyOrHNbm2PpJgBQR041LEEhFPS4fhDymXSgvr7HAOKRZgqkQjnrn3
44CTg58oyErUyfGiVX8Td9CxqNsdSRIWQ7fv6QXRQ4IG2g4qGCPfqhG7dpbTTIkcA0jtu5YnEUB0
dFIbf8y298ivjT/TDH8JEmT3cmNY+Sj/S91+bhjPZBRKEibNubLY6PAABlmB+EVno0gMHPc5g8KN
u+tlZsfmxHrn46NmVrx/TDDIH9jkNza+5j9PXqVWJFd0c4qb5wdMfTiaAfjuW9zGYLmZy9pPEkgQ
8MLbFexyOH1TO2q4A0+CXqiq+8VR86DIPScT5vquECZBC/Aip6hlOLHvjPuxsz3+MLOVi7ukj0WH
N3gM7d6OmVSvDqSxuoqFJ934CYO+zE9rjyRYhjQNMFczJeDkssAGhB+9EtcyrhZ9EsGiFmuqJ9Oo
Z/X6qWcpfqvGIvzCYIFm6VXDCd/Xfdr1Bx3VRDwCFeiZFyjnrMlznCi4hxUblrCnaO6M0gPNZRLS
GBQ1BvuOfoF5xgFuU4yIi8skYJZPTnunaP5jWwTj1lbCNEjHFNP4RX9fc+pQI3H9kkkB4lMa+ll/
zyftVSflA4kgjLSHho5SNVyt2aomgqTywgavppF9EVSL3O4SCqnGB7P6Hn3Z0BDaztO47Xc5DEDk
J8yOnTp91OwEg8V1223bCoed7ZZH24TOlzDtiyyuNyKCbZQnSU8t6oS3VQWAnZzhaxIkPtdSUsgV
ZTjhPYD0dCNS+c7OsJ52qKetyAG1asF5MAOz7VGX2VtzkZM/jpXOri3DG6p6ygMetiFKhX110FW+
ZtRRTeoRvdB3kmNkkdJuy9echCZ8n9VQ4ZtGmPXexH1N4YRidv+s5SF6BF4aD/y7ocNmlHdH3548
pRkM0QC5FiIKYxLXKZZDexl0EHy+UZwsSVDb3RtzepHnncUDfqOtnoSTMDwZ6+ogj2lgNpSlvu1E
YALXDK4HRmsqXnMIZIJp4DkS66C/GCLMKw4mo2YgSyEwRuQBRhBEstXEOAoN3+jq58GS7umHd+8I
PNf32APO65B+dsaZtkRTUg4oV99ZvVvtZv7XWsJKEqRk61VzYF56Y/3wIOULdRBms6gIQhM0cA6p
sRnOop/q1yHiyvC+x3SSnWT+A66WeXXZT4vCtIf1SDpBNCESphWpssqI4uuxZyRQLcwPKjZ2nCnd
ZJ+NEQSpOppBtWc6928F7yQcB22pyWCu8ALxjwhM74Uv+HINQZTV2uRa036JPsVsCv6oZh9zFbeV
tk4n0qsdIeUxUTRUCu42gZ76HQN1rkDHqsXYqVDl8XwAh5pCJmdYMIWRbvIp2skEfztgTWdJF/43
W8NRHtor2l48gD3AviKFaS1Z72A6v1d7HdgJvDtztpLvO+y3X1Wrb4M7mcqJh6udMTJVHHCpzwcC
WrW/PFG41Oni2ixIKc0iv2Uvpbz7GuMSCSaARry5gCDPCZcplPAsdOm2+eVzpz9+f04rF/l86nQA
kNdM9AeHrs+LJJkvEOfAmzqx0JaU4Wn12ZiqtmsPMkpHZ4ZLQ8VBaaIRt1u//Nkqxt6krUJMUjPp
Yr6V50qnGQbn5cH8WYKAkgYhsSpQyTqJEjfQRmRW+1wZq94FCZGWYmF75mod1kvIqsXy1DS9tf2s
RBCMqpNuwjfcwCd8umXtFjQknBxaSwm/h9Zknk6JTOHwcOc6AJxTtaMfotl+EVaVlAZn1Gwu8Qtg
BN9tGig7OakJBnW1iBEPU86wUP24oF6JW8z4wQfUP7pN210APli4L2wXSV9pxby2W0B8X9DKInM9
YPAeAI2zNovUEFItw0KU0KQ/7xxc67kJzrfrkrjc4wurA6An/Qagi3QOi3xWtH5qTFFvGxxU94Cq
xqXQIAAW+YxXXNr/k/UWqC6p5Ys5q94c5spcV2Xu0fkWhjAGSCffjR+dNKbW84OVHhbgT8+PTHM2
z4kMtWA15Pyk3aPoUTppWtAS5/oEYVP1yGltCAkI5UC0UiooU2vDJGC3qN9v8UK1bGJyhtQUQCxh
zJGfP4w3NR6HkXj1i7hdxmGufvDMbNW8nt0FjbmOv2XsKGupix4CB+LqgohjQYjx43eD7+JiXGyc
/LOhgnC7JJZBq3bp+F0SLAwEjeskOx8oPcmXIyFB2tVwQ+UjfOIVvkGGxUnQQJ8C4Ar8G0S0GiHB
OKp+8fEZQQGU8OocmXU/oBxAgmUtKdkj9MCNA/e+MRr4QwQPRS/xwQHcluNl/jUcwxm2cqIF7vNt
jJK9rcW7vpjNBM4ZpUCd7wBxUJUXnS5dNmuak4XIdhPaikE5l1UcJz6JKkJ3WudgHGpsFFZ4o+sj
wgsRYXekEaDmD+6/ymDtvSOzwSEtajVU6G4Cbk2QiXhI+cewVr2c3RjtUjfJqvgftr0mgXTwiCQU
F+6PP2cbwJJM5WJnLyJwLHglleqbHxQd8WPlE7ln5hZcxs5ZpvZvfD/hOjcBbd7+HBbHulZ/QIlX
sA7cza6eUEj6mzq75nwTE4kw1/omy1/KWcfswz1CCLUKezaCLwaUEd6ApVSNMGO+nHcGIA53DLBp
33uhnMZPRnM3rGA7DvDV/4tw8YoldEXPonivgsakmOzntHaZA1zTtXSbSd/NzFVnUyM6ZuzxWgqV
F27ko3peFqVCzMge+FedxLFg2i8urFlJ0H4fc86gw1YxFZumCVZeJ28yBKQ44zkcKWxykqulgduN
AZesefy3DPEIOyJjl0LRbrbQ37j+0Hr2a2Wn75tIjFKU90ErGxbEot+kE9/C0rSbglp5IitNxOen
+5n9uCpM/9tMveAqOAkefUCh5BTJmfJmeza+9bgIR7vKcpBDP2PNGZnCBGgscl0ZSEC/hqwlEXhW
V2DASqil6OIWcFhTfRmExIUNGMAInR3jX1p2zqZ/imI6H8Qmo4za9ERNnWq03Uu7sVFFdOGUd2Gl
08wYrg7fzrFkvRcjyGLGI7INhcDqpjyzXraysfv1YryaOPQlRHGQVa4CraeFaM/LnXzT2ygkpIXa
vXmtwRkfDjzyDgrZgAvbYToOyKW1bkGy1LtU6i71rSEFRdON/AOq2oG/DsQyn0fYi2TfJDGOxi39
kfbCz+fR5aDwn6IK3w4g+05txmpa/8rr61KNr23KCO/qF1kMK/yiCqCMnisqZWqdZpBJjNZNW828
D/vssC/sbh3GfCjfQBcx4ZRRtCF5lyJC+eX2KiQIsXpUQCsg8Jq+GJ0xSE3XKC2JvgYEzvCNR2FX
NSba8FrAY3vaPudOgjypw4SCSJVqjIgFo0jE3rH600Nn/6425wCQV4qGUQR6zcruKljXJd+Znwnb
xUMWKZfg2CemNtNEhAwcCb8q10M0PP1ulyteNtlIxWd+5peTW8M+oCsJGF73d3iTkNAHQuCyxQ5g
/0PauNQpVZKkp48Kgkr+kxP7U6rpD/QQFgQhQTGmktjvrY+6NZ6ReTJlIRjp+pKA9PI9lwoeEw+T
l0CgX80IW8H0/09uCriDJod63FLLHm47SWodv/6ag4SkER4THF+Wd3Cyeb/8hV39DVHU2zr2Ft4F
4/D4VmaOYzgQhVwGFOBeWJmwQwQ2unuF8w3tcvgUfqtWFKClVTXq/HJAVJH1YTMLDcja40NmNMF/
4R0R+eAUzY7TWneRYhqWISi76R+UOl5SFGmWxeiqwUQb7mUQlSobzWepmvCQd6NjN6Ew/IEvsZxo
bUTFmi3av7E+VIzhoqq0ViEDXz8PALcB30+exJM3Gxpn/w84fPfjhWoiKLRbyXLEcd5VUNBYfkRQ
h4WFcE45MAmk1tz15JhrLH9gZei6W50/YRhluYnOupF+yBZtg2N8GRV/MZk/k3tldv5UM6kxhTGG
OP2/DhFGqpPFE+ZFE5IxgEfztFV+CFgD7IMEaY7/psc6U31WXjn/faysbLhBSUMCVE8CfM4QxBH4
TMAaCnheEKJsH9GMGHJyMxR5N2tXGYhdQTL4C9gKqXcdxDqcqrbUvLnRA40OCRMyMKCgExKNZuwl
SwYQwzqwH4AQR1soZB85vLIE5VNLEQvQw8ZgF1oS0/2i/H3anmEXKZGVY/O6aN4IS6iUymegNFm4
l2tvbUB8QuUv6rLYnw5ZYwe+KN+IDNmzjYPiXZ+57KUZQVSRvFZhKVyDk8HmIB2W+FP6G+5JZO6l
YJ1iUNJFoAg9SoLcB+kW8Xs1W22nb570zg8hd+pGn/ELDSSMa5S+llzx/o2Cxp5+YyYFmsNJNtZW
T/1kqqgFsEk22P8dqY3JMEpDCRzozvq12NRcmVfUcE6teTtg6IJTB/ScgYUhgK5SRQkmNDdKEqtp
FUm/HhbRav/sTD406IkRj59Z34RyWSjKXbHH2C9u7XrXia+BKMm+p+WtGxeRrcpG75LbyCyVnKLY
8aE9S4M+ayNks3ERf6KhxoqY3FC5+/r3qpsbszUCsdinLMNq68lBC2353l0YU5/wDli1d0YZpvgM
s9u9miVhnBdzQqmYx56yBhpPungfcoVlDX3m/PDa2EV6smt+W08Z7JcYqc75UP9OmwECgw++jWgH
3EQa2sFTq6fa4Riri522hCqOp4h6iDt8okr8WJdm4cagdkbAZit1MF2X9XvPV90m0uWX4iT8SGc9
mPgMR2zkOTqAL3mm0RZaBAcBe8vZ1D7tPkW/SLX4ucancgR900LGZuzc2mSp7X41MESBtOsYwqgI
gmeX8y9pIVYTMbFYzXNfSSQn8IFRfbCCWjP2CdSVZb534W8u3epMU6+Ags5evhwLFFaOpFNaz/6M
IM6qL57toDTBoAUMu+0g+Ct7BsOHbCcfCqBPBb/QA5XRXfJMcBlAqEvrm1ctCuljxLmUbe2C4tbw
OsLda2xyb8+VRvRjYPZb+zsoTPJuwf3kUQxEPnn/HG7QZxiH2TlaKaPj+EfF/0bCNLBUObxgWpFQ
5PENNeSczxDEkutBwpNW8nYRNOUouCeiygYTCHdnI76RByYIvDXobdTblG+G08YmrTrQP5/cJFjx
in4xgR1FviYWToL4FG8uWp2breVgcRvUVvOalRrfLNDDMLZvZpEmlKr2rSWiOFKenmhbqyW+t7j1
arjwwBxZ6YJtmgvQH1md6USEC5U4oshMwdjWKEzwC3xChrDXP912c0vrqknsVKzLoBKTYrB2qMZV
Sw0JWCvBvooPS07CW+EXs5uswZHMgLTLpHB/Ner7Ywtd/VpNgoVmg5NkNTVIwVG/srHE0ljBC6EZ
aliy6gYVZLKLGJsTi5h3KCplmsl1SXFvkRtYDcpYlRw1tTFGpcF9RLpDTWidF+NGVYlLSgX/HHTr
f6lh8CU5Qpac0QK2MpgIs/0METyt7RTxyXuDdozR6cPywmxQg8RFkQ55wII1Yg1844hOIW8OmCN3
1TrU9cSP742XE53HcG+i336ELmOAsTP9m2/gYltMt8KA8WfQuCCGzO04+b9aS3IUFC5wLROui5T+
BVHgVJOZ961Cc6Sr+i5meAYHZeLLafHGf5OcTFSCm+A/+v5CKS9bxzUzj+INxfs6cFqgS/98q6Hw
Tk2uM3XUDxeIs3VEGA80Vf+TCTZBZNsXOiQ8lpeAcCXTedmkyY8+kxGk7/THrf+6jUldCD0kkIfX
ksMLMBd5ZERlOk/vLBz3o0t59FarLesZVGg+6KgcSubJ/qwqYoLI2MsSi+GFe5zfRujRKhMU6NAA
QItzLBieQlSFP9JqxbkuS57XdpycA+xSETNzY1oOcEy+1mauu0DqNtwdfNXmmsvKRPRUxpffxoji
BvXBlxn6TYvlI5whmhWkP4iAPW8ev3do6jKjdU+Td68BQHvSpPOuMBcybXFR4X78+m1yqnEPGghm
FJTiKnDBeiilJO7t/ExOPqq0ONNLN7iX6aa3VULXAz4dJYdZJ++l7FuFUQQYXd62UkU7PD5O+b7d
LQW/mj6AC6dtxKJFIJqRO2ZBXNkgLxZPMlUfixk2NDkyMAIWllXgy+AzE1kMPFV9S60l0sId6p8F
vi/bx3OnIJNU8rLcN4QX7z+c/RM8JUWRmNYQLaJoQW1NvCcxN3nHXMLQHeHxdA0lObbz5AB0Ju0X
OJam3a+odGsNVKqyFN8xgx9gV2U9s05+L7Bo2nw4P+uNKmcjtvPjlrxyd5kNqH/NppvQ3w/mtxew
SaXEZnoNW1v1kr8gtcynYUk8xJlQd4WDZTPEUKk3zXPgwDDpr3x5SRwIxOvrb922PxHPLqlSdaU6
lZUikHqpqtmPTz20N/BOIyOSSYmQt3xUJ+m1PfKAni8YRLD1UkFCHne9CWpw0KWm/fodzHzeEPUP
w1SIQJIoAmmwEzIPpU365ZrXPhmUqXHo8qTsM6GRWMXLcNAobGu1TWn3cIBEod+ayaJSCeVJgKaK
CbIY6NgH1GQos0r306M+SSDvRr1Ihp6SjKF8Bw248MLmZwPtgfCv0Eh1wT9JKhISL228Z42npr0C
iqRYeWusSDBgrEdZA2rof6HMqK53Nc0RysowlNR+VFUwoQ93nEyPthsal4HV+gjQSpsZ+jsuoMtn
gDOb54akAj5/VzpDy+qwm37QFquoBWPlcq1ftlRevwHArAD2+NoUU+/QoMddKmYcdvSBeode/b+3
vMSAQih5rzjI8On1+uayDk3sJN/O6IYJcsByaQ8aXpOre6moT/0GGw8OXf3vbjQkp/twiHEkwE62
6X3a7gOqyvN48+Fz3FIqoeux9NWQMnAClzIBrd/94tAbGmD5HuP6+mI/LSSK5gRzD91XjRolUIqt
lQmsGop8Mnub3bVhCeTBFdOHiZ9EZ9BgASCL5ErY7OgpOzpBd+AEurEBcmqCjXXoq+UAvLX0Di1U
ljw2hoaS/PneA6bmetIsdmA776PQqMXF8BKK3ggo3JH4C0eVV36OUmtTDUug7bHG6/WfIdJJg4rZ
6ahTNT+b/FObc5YfIFvR2sZKNPfrITimU9LkDpHNXEGOKymiUibqmV+K58dy75dPHxKe/5Lix/qs
PVTTcavNjEYZ2eirySJSKLI78tMqABMjXcgfJT6kwR4uSn6/Uv5PXxbkTHYU/I14zjPjHoWjFyB+
AUYio1ahLmncMqPYwmBlJDWm0E2Ww70VNc+LTxs2Rv5pVSdGO00wZKb7NtTnxx7kwHAdRqHZT8+4
PKdZuOdxrcjr0uWrrcEi6WuZ5+uNUSV6d7vrd8X0iBd41gQR+nEwG6QFRteHXLwRgqi/DgUezQiL
joY4RVAtjSmmzhG7diGLVb9HtMiAJLPUDe9r8iHIO+auTrhbvwm8/bzmKXs1lLhFUBJp3wvtsZ14
Lo+qU4WH2vPdiNxZJrXy+P+opgs0VlnNerNxOU7J1fYUf4kQ5yrR+Uq8Gg+xP3HmHX8xt3lbggI/
N7brdGEruVwee2J3SavmZi168QL099oF8pZSbSEyLLkCBzci20iThwKOt9Tx3jMxU7Riq6sy+GIE
X0cQ0lL1tFaz8cQKr+1yzad9lDoiA7PjHlRzThejozzjx+13dpf1kFdcIm9/avgfKXY+Af8jX/oC
ruRltGKeNk33n0yptnCqKa9mKs62qDUquj+D+pdzVgT+L0Dyfm+FiV7vjVi5pGuwhXMLTePgXJ3j
wEV+0c8fJaU5P5D0JQrqqaTEsLf6tob6cIY7ekIRaGS6VqwiaeSDsxyb+AxEEU8+Qge2uiQsbMWR
4/gZoE1n0vTLcxlEqmWnKme0a31moT9QTgxF9S/rYgiKQ+MGuU/AfFt8iNcScTT4BmD1wHIna8xI
wCYjbD8huXHgNQJL5E+9QEwB8Vtg8Gj0pN6ADt/yzQGHOHKP3RZCBfgLafKzMK6T1k385Tjqt6iN
hKDXo5bK1lm+kPsSpuH+dAXZEG9kMZFZZFOpX65IoWF5HcY+zyoeLzYAjD7lsAXXOkuWkEiqxvIw
a9BUTbZeUn3C7qo9wf7Eudis5rH8Xx9LYLLjJNv7jOCyVVHamImVXo7X+u6XLjViarBRp3lzq7kF
yxxqArn4wGY/nDr5xPRXWCj1O1HkmKmZ59KPYZNrFw+z2WQtOKkWpRBTEtdZ5pqdnFZHX2zEZF/R
ZHR8jIFmINmmEAomJzdVX6a8RELnpOHxs6EkCCUWfMIvcKbttOxQq6Q5QzI6uHGcKI8UAou5gRO5
VvwdpvhnNeQtvAF0MBOCt0SN3O9h+HdGqekcJg5R7fGUD8JCniYCPtiL7w92Whr7H8+TUx6MjR2Z
ZLNrSRKtPvUU96RbGMWyBdJpmdo+damLdw9hkzkuYcAQo7JdlcbsMdMNNRfIydtyfaTJZfzfFDcD
nStwF5ikoD5NwnOlKvG4J1RmG6vzLvxpHDfqBYcl4+ovGQtzI7ad5hiEhMeRxigI99HjG9EmS+xa
tqurmsjIeEBg2QT+2mW+nTRt4sQPjdeyHp+jpDYU6VgEYqr1VqVOjU5/REJfveG7TGJGwyDqlNRq
5HLVdwnUBPDNBEFEl98wTuqB7j6pSFu8k24ssMK0nMnUU60IziNNhaGzl3eceMBPTluHAHLWDwXN
sGorG1tm+xFFJUc/GV08RFGYp8xenak1dX/ggK3NSl/TWjrX9jl1/IaES7efhi1jOnMIb44S6TTD
nMNAqQtluzleVgEPE0M0Fwnk0gO5L7K7Xm2/xdmZNcAihItBEcgiMFW31b4UB8fhmEbAyaOpG5oP
GJ8NYdycVetUdH8t9awDTy+4chMd6ZjAe6A6J0RB9Vyv+g2rbQ7I88e5jPwhggtLHVlbTV+60/Sd
nuqax+noZ9ECTSQtdLDzOBQuxRHexsy8ITCoxGpEIzRR21/v14z5ioYGDcCd+8V4JWEFINMNiMTK
z1cV+jEoY5SOvb7snoNrn22QP2EUq6PB3WUrejtVoGU1CDZTthuIpPTjWYBCw4Ip1XSNqlx7eR2F
JZEc3d2aTudIryjOXAqob8bCFKfD89XE0N1WDuuxIatov2mYZaap+Py/RVUc49MyU0XAnE0VDeq7
iOxo4PsQBIzSJR6cf5AdbhYxwDuBpwcT7hUBqawFAAtqbtc4K1aCpqfa6yacXuMqPs4dLhNIhrQK
cyO3/n3u/Pdg+bVg7X00LBFW7wvaxGYeXad/NB7URPb5rtLdWFAv4efiM/wscS8BrnS4wSdaSBCx
tMSER7IPIw3aaKGTntV3+25M7qz/RPSHBC53vCg3JKOEzHJDSRMGl0dy/ZJvsdODx+6zPjeZ+p8M
ph9XY4oUcbk7YNfuAZD+XodBVzHTX7jjwddkmmaJ8XuljTUr5/fWzQRaTGjOBwugsTp372JwAIuP
ckLV/4HXv7x12XV6boF7zFYSdn4+5agYMaOc700/nb2fWueGl6fRzSgtKILhp5Wt3+9l39eI4Txd
/5vCruHaDKTYGt1T+t3NhEUy1h1xSULImvlQUNHleQezTC4bLWwvM7b01vYhJAYhXRe1T40NruTC
5a4q5DclUZgClkWtgStra5PzoSi4/BPI7tNQVmiwXfRPI8fUD3OswX227n5aMmFQtHOQ7Pbosshi
YgjZ+JegbFoifbQXmcb/J9y7rEe+fUHJcjb3vRpV3o+nNVoysl6ZhXONufnwMnlBxPDBXlpbj3F0
g4vhPC8W/vgfQhM2GoSXanXHpps9HOQSR1MpIiv1ymQrWxyUyFfnozfWfGjI6sCLcIdDt4jjLUI4
QibJ4ytdnrJPuTnbO9FXS/xdIcqqxcBn9KyDKItPL5/mss/RQG1E7MbbOfXhCd2eddBg/v/AwXE9
77QDXeu9nz2pc2c1fvdb7dfCmucH8qTw8ZOxQSXLg4yiBVBHgM4AAOpSKT+beazGkSs1Sz5xxzul
xSAjAYk0FCzH0aAxm7vo2n6NBGODWP0EzhXrLRlAzCeBfURGXy6UAqLk3sFyzXDw3VYi7Os0lcPa
n12JDVo7KCnFyXlAmk+N+aeA6RynQX1Zwj4OHO3kK1q4SF3CYlIVcn4kGCTN5fun3sJYqTXjBPmD
1J5hrWMnyVY4kIDYYZmdR3SLP9Xlj/G7tvJaM0rOE30ARQUwbLtDGjH8jDTNlDbp3MPTOgjxqa/j
R0KTMyeYDfQpa5n2kCrdY/wEecJ7Pix1PNrJZPcYp3gjiV27/fiYA/RKu6/y/jlNljzcvE6+rYx2
UhtlVuJFUuso+S+/cqvQIMBdt+EBpPe1v0Ze5aI3wFkPSpdgtoHpsb7j9zEUNXvNmkKQq/blyxSk
JMrjmNV5MDQ2HIx81SVqok/jWdXfG7Ct8/HTDTu1DCdum/T03hI4tfLHKzN/CZytCqXjKeFUi6KQ
KSC/ELiisvGhLFg5vyPENq9FmKO/KczrlTrZ2vUIxAqsFiKBqlM08ynNkla6RpGRc1kdnxiOx1C/
C0vcbxD6QTq946JNs4X/LB5yde5R1Zv5Tp6fEeQlrwkgL07/v3w7E9LBhjv+WPTwGbATQDzwjpCd
/zGlGV/43DuhhxL5HZCWo3XzBT7yCKEbS/G4XPJGurruXE9ZOHJ8RBNetjJMH5mCE/k84MEJO+F9
lE8jSstc0RlAqw0DkIOBAIZ3Vtuu1H6UxOa+aVSrcEJMYHGKmzYCsosPlClPqovlm1dMBPa67EMw
8H4BHbn1ec0951iSPl9MpXfUcyQzHMTKcUHlPEEEecpF3OBQ/z2utJ9I+fTHJEm+PBTZsFTQEtr+
bFMRmcuoyZG81YBDX5alCL5FWxXWlkQzqZ0eXD5DMoJaHYgom4dStmwwXqJtf0cpZyZJhf8n5RRn
HYHZCscIIp8Bw+X+PRb6srMRJJHE4FXhmoVQHfJCuaP/0T/A41b64ADZN4DU2d4RqT/oV83LW7D/
FYY9nWEb4vhxpwuUHn25+fSYP3hoM2CNRXSavv2Z3c04pMQbQFOX5PILaumBngQ1+D+r1X7QgRlu
oFZpvlVoBx3FfkCZbxLJ0NQ69Z2vNQ2yDA6PLyDl+4Xm/hpEIrntQ8eMnj1N/l9QdaIigoT7KW5B
FUct2UXvQSMvg5Ie+wSu7j6CnX16ybT6KHxLByfynXr0AVIHbw6xf1ZOSF4HF5RrwVrVf4e2Warc
vzTMiBt9sLzpP6cZv2Xc1klhvM7BGK8AxOYWEx/veKERPaz7hacBKc04xdYEB+0torhCZTHy0JFA
LwjlQs1gF5p5Wz4UirLdKKCIkq7L37EDih021YEasM6VKOuFFOosiIxTz8Mr2Nyn+tTLbPUdBmpy
Kj6DNUN8aKDWVenP4JkXw42iPH9vkD4PHja+Qv3IUmxVt6GYjvnysEckZIH7G+M8JHMNektKmQ6f
ZAm4+kkjc5y4ePazJzPfQNZf8hNDRFZqiNE186iYyA8eT4fQxHxoWh5wWcSBrbo3oWgQo0PGXORO
spxekIweO0FS8NrOzv0tBxSeurH9932hmHmt2e83ePwCI9QOMLxHP+RyXCm4WqPtDdSZEks5Obfj
XdUbr7x2La6gaD2SocoDmGKhQ6KtyUsKJSaM+cviILXJdXG5sSySpbF03aCJYNtOCJgQuU5sVtNj
QGjpqUQuw7oxpD9X8C17yWj1l+/R/wKCYdZ/qZ0S6iiAOGGLyjk2gQDbAM6/JegEvcU0x2U+yHYH
CQwMR8UAQut3sgDx7dGFST9wJwC+X+wSPXyIJvLxCG90bABpU1s0fQxwFxyqQq8AxPxYX8X3qvJE
+kqS9ekngi0wdl81Kv4g/yieTNjntcdcRnumfY8GdXVoEnrtMIK9F2+S1LboGzBVQ60YMb2Z6k5G
nU3nr19gCwb8WnUR8VORH2CXUjCisVwtILa9CSIdyiR8AXirgWdgqK1ikOTrkE+Um1P0VI50NmrH
U8xPLwrTb1DLrQuxJJWTFKapl75TaxRlbAp/1wBxHd6zpOrvAOM8dEjYdzJ8IET7godFItItSG2u
9WKfoK96DH1E9ii+J71bb63mKUDqc69uOptthk4PjzdyPk1Fa0SjpvR1nE8yy2A/uEUMY4NoaWFv
6TOCaKg4LzndTjns0d62BXTi2egMdkWaJ6yfLq6jiSU6W/54Mk7YYdReE06JHgt5xDtkfHNwwJ3R
H3i+GlYpWtKpRkaQj/f6Iw+Q1Jb/2RVKAQytekqgrmZk81zQpKvpikqBTb4Begm0qT2pfmh9ugjt
VthTVx5+UJZBd4tb2NDrSmp21l6sdf7wtMJqiWI/ag85su3fUbUgtQ41MRwTDJRlQMy+pWxCcABb
60rbtDePm2ZRFXiVkGn3YE4zMfr4RNqSnAuFFDXD0tfu5GKzu390AOFloOXdjp4RvWtjpeuT9v1e
DWQb8pKQzJujTiqRmeLlXtSIxKpaQNRgU+WQ111wANdSA1VzOeDHe+/V4vgRad9m+z4qhpMhOSgx
1y+qG9T+gXNXjKrogw9eQHbhKgOjfls/QLYgc70t3Q93dYicwWFQeX98mfXSbU8ywzEgoDnKI+2j
ZSja9eTcGtIKYQETreud6eezfaTh4+J/4Z501e87NrTQoHbQRzI2sWMh1QsYU/fKQiS8InBbMdGW
tBm10Fu1W1OUP1Fol4lRy96WnQPaou9jlOV8q1stQPmGpE/5ziKGGpo+3De6VcXlYieFUkK8wnxa
2DID2YhVUC5EiKdjlXdp1CjSrDwf+7TryJ4P8RzP9R3R4Gg70+wYVWMFYl5SV04iwbfPQJ136YUQ
nFEncKgMbr4j3wtsE7LglKcLqLuZq4PkcRGN0OwvfS+kN7kHbPOQvAYZeoK/aVbjkKgmwTTWM49E
KbJq2mRGmUVIT3HaDBnFMht2YR/8koUJkZ47EfzKTbQVIuxxMEYTEVfeiuWRjC1539ybW1MDIBL8
zaZkX5wQFA6g7ljG5ZAw+nmCctInct71mJpPacjmh/FKE5bVj5dK8e/k6Y2O7oDB3hr8TXlQ2krn
IBM+pJ7axEsTw8SOU7c8z4fqG/gh1oKXoK2niVGutPDmSUHkN71y5K1taGaSe1EXRHMl7Lh/Wc7C
CAQ4uRzDNscZUiSHyYTvNAHImSjDVfcPhsd5n1IL98187v4cDgizctN5JPzDlHKNTwHTGXF2HLK2
nWY4k7mzpJLtr2TUKgnZkersrTI778LYP2uju6QIXK/9F6sn8mE5eAmo9POze8+jCqj+awu5ngO0
2I7pQwBcMO4xdNcHwQ7kf3+M4oACPyLdOA11S74jxFJydAcK0alN+UU2wC23Y37BSI7hI0NJ0Siy
uEPTOV4Sr8RtXinStUGTkLxu9y186cmRa4fUvcJOLRykZ0D9SM15vqawfc66ZwS+T63OqMlnuaPC
OsyDZsqwj4FU9k8A9nGf3CwnWIaw5heZzffjqB5iEBEcx//NO6okbQk4GltDoccEgwitUIzr8If9
PjmJBFO6G3GE+lYwWYpydp1WbiMl5RWFKyy/nCckrDBNiGdeUoQFZMrFc5WgjecQBZv8HhJKqVXY
QYHAzZiUXLGeKATuwpGkYVQFdFXp2pjx8QIduRAzjlTGadMqAQuyejD6+4AEeoOHfQNa6s37Nrks
c2fN7mNx7JUU5pqlxdbFlNRLXHUgr0DyoizpVqxT21jgmtGJz8T4Trz+L0vWJ6vhiIxoiyocwP27
0lTTOjhSwRuXNB3/ov36YV7YdqWzfbuYiS0T02QhZmYjsYRSijJY4iTkjnNoqf8XW1gAO2SuYXje
VMPXsWypy35kqpKr11zZb/NUlv1K4eP6aqIta8vWCJp2yHxKqe82BFHGXhRtipBEooNUJSVIBalF
izY/Y0/MzlzOzizG5V2eEWhqIXbr2hZaGHtqEMqLk01Oi/Tz9M/DmS8jXD13d5g6yGfNO9PWcogn
hXst1IBvtUE3wkqONBBKOd4YNDchukl+eHiTDuYpNmSP0B5/bcJgzZkkKmGAmYuKVs2YN31G3Z/O
aImTnkQPFwKxR1EebCdDUpytaRKDBlOlKDyjbrdO3kHDQ8BqBc9aYRN9fEPY+e72z3UWKV9S2oi+
EfO6n99WM+l97p3IshepILGxum6YaQCDEpLlduNtD85Ba93dnnlL1gnES0Px9V3q6E049aYeBj2c
528Jq8EUTatf8CVdBxpt21SEVs1sbOw92XeGxZMxcDd3ecWSKt8YQFUtTnT62/LJ+EhovQaGeR/t
eE/6No8CfhxdMRy+zKt/ZKjuCyXse1DB35N2iiZDDHFMd4wUCkLw6NtVxCmVlVbybPwYks2tfWb4
7ogl+IGZNDylxOTa2tdbttFXm9z94DmMh9NQl+ljS/3vsX5KmlyVBJl3bL8UzZqxKrOOn2/3pfmv
3MaTeBtWok63SjE9JeHVnuGzkzaI5SzLHmfChmOiEBhLSWVtjdfoJFpXxDUGgGu8oPIWQD0YOIPi
Jzre+AfHjRz4R3ndtqPdHcArhh5FKG6c5Gibnu46ArmSmowIYcKiSSe/RBkjpMQ6JZ9E4149Rt5E
hMsFGWh/0K05uM6eGnm2AFAfwvXe2jpcDvwxjmvZeSEitd/neIanSbwaAbojbc21tWJ9M058G58v
FxC0Ql58wmuOJSY2nf4j/XNVobiFbX9qHOB0sQsM3vay6ad46DbCyur8GCDyXIzE0wDGFDTX9Aut
ig1fk4ifZx1PnPNh3jV0Ef9dXdfMaxLNulk2XZLeTBU+hQj1tTVrQ0ElwW5G8mb6iVI+s7PauaNp
lx+DQV3d1SICMFd2NraYQXfZyWnBYlOFIGMYP1PLgqdzKpPmooWZTuuRbvIvLqWj3xep8yCAdg63
TNh926ckeMmoT0y6ozSx/HAq6fUhTNH2YwCaSGaTAcYQaDfonz/Bf7arKjLjadhHdbNPJcSp9ucS
40xaRUp18D5A8s7aCIp8qV+okoRBxT6X+UpZmQcBM0uW3dSTJfr4RCxl0hHy5S37GAb7IuLeId3j
Dll03JYhIuY77x7Aje8ZfGkzV/HB5a1KAYOEPTP67kQO9Fn9qaJ+JB1/NGtF6dL4pcsuEQ9c+o2e
dfNxc+9KiMQwaa3vwuqlWEw5xMhSlzbUsa4jr3huf+W7cfTyF0gH0yufCC2z+K9/h98IQ2EIUwqv
d2nqgyM9fF1OHlM/3LMRZQLB+YwrmsX6SitSNP6/hKYnDRm8ZgNOCC3hDsp6azu5JODc5B8r6D9U
NVUsnH7/lP6Xy70sjWphjeG+MLJ80dzr8ntqXiTbqbsEjv8TohM8JHDOV5dGiNySv1VmHfylF7I1
zCMN33I1tbTLHQrNir1uARqCE324kynjRd791d8eeI/yyYbgWKlPvbhzdhrV/okcgpUUb90fl8PH
yNH8nFmPA395ul04pRF2wnfNj4nxkobGZAbiXaOlYs2UYeNSTvbe36BClic4EHKJlnW3HR4vfbSp
9wSwOfT+zDsfuO7HwEBBHZ3iDeSpqq1VoZoLXnYre3TpuA4n1xFj+7pHHNtbhbWk383RzEkefxNM
YyJU16w28+Yk9NPhF2EEs1659dtKnXuS9VcQVm7baYLz2yLq7DJvMe38jnE5WRbXr0etOCmC7V3d
hqLbHTsDFEp43Pl4AWExsjXTskaYEcnFcUZePvBoCeUjC9AQR2tmh5yBV5LIj2xwqjcG0fFaiCCN
qxs5mwIYIdpCFRRrkR+CEAR9nUvwLexFlMhNZeDMHS4ru8Y2fY0DIp1DqSJnwXsW/yXjCf90B76z
Jo7XvNO2KkYruc8icUYMgAJQonJgkolKWxjtVn61/MggybZNeu3lUvtVwqnYiy6NrUW6a2hwyIzS
HlbjHXHSqH40w8EGsghTeNS93zTn0hSmBFiWWD564gfUnQzcRH4IPI0+ghrLmCjneUsyGsgzRL+9
q07QojHERBYX6rRf1EZ6hGEQOQihBf894D2qllxe6j+rUWKGj6O3NSNZSVGZrfNIipf8WNcn9lse
3RWQRmBSMUPyBkxMl/wqffc6dHjA5gOdnzGgN5W3mJCeV6qAhFxMnirbbY7AndHYvsE2dW8pHaT5
JhPPNFcPydzWg5xccSejZpU+F0mdBuSz3Sstiiuw2XQoBj85dVtqpMoWAzW887G13T4SEwArt6yj
1UeV9QYaEQ+4H2xMAq7M8KhBRNnxjF4Dnr79KI7iPMJMg0jmpHIwvGcpJiEVHT0hxUiqm8Iu+i8X
kx1eW/NhOWIk41RM7n6p+xDboxZcCW3qvs4ogVsosu/x8xyF43iYhqTD6QgSlRji80L91b1YBq/H
ovmDbqfpVmZ4sR/Og/wP1B5T0FVZLRykzCaufgFKuNEPXoSAXCK/ahHRaIoRQkNytLqbT2eMw/wl
HZjc9DZAf9e3A+KoCyAWqAjV8dQjSwYG5WYhKpdZG4xOqQdyEjjzCat8g5IzuhcrTDHNpYcPBgJo
4BTNrGYbsWtIYcaQNeFuVUmbVf9jIL+YF0dwdSM7JYp4lG5qapYkpat9ttxitaKbmFOy3QgusSCd
W+d8GZxSEliqeTGk9vyPrjMwTcjJS8QynR+Qd5pEIGwTZGTBFOiGq/Mk0fZQnVK23MkF86r5FMAH
sURQTA7126B2lrM4yQJEXNLC4o+i8M3NkSwLXkW/jWwqBdtIK9C+MHssWdcW21pikAzIL/i/Ua+P
gZ0enAe5B0TteDOOT2ThzmaZ/AoDIQey8vcAY8Uwa43pHvMm9uHl8iV1ZPoySG8FRoH/hfrPaO0V
bZQMB9CpRwaP6uj7MvEG+jpmkLmUqUpJPJAZwOL7icM0qVqthGDEZYIo9Pxt7SvSa/BGDjZzco+D
6tfEgUaytIK9DxDkhEB3hYyOwuNtrJtv9I0jtrhzhDE2W9dWpsh1h2WB9wJee+LmFkpxn0b9OnyS
0sd1IeUTO00chcTL3JPpvu62Ro2UB6mapfbw2KQqKwicRs62c/wVKtiNBFMz2yr5zJr+CfSbhjst
yrcZL/2oty9q0p90a5CRmC9XiNf4+la/UqYBm+LCiKXRsnzgRjc+r9Jw+wBBJfHTB5h0nbDpJsd4
33VTN35FJtj/V2fi4B3bNfHRaYXr6gzO4HA5fTbN+MCnVyt8rCJa4EnzFiwRiq8gd/NbiKN3HpxX
Sx4Tb4nNqIXo8G11XYuZXXZScw/B648SVFV1ppWoK7t8cbNbwUagpFxR2BJx48IRHUdkrWR1Ze+b
B2BdUksrcJZjRbWhb2dpMLPhqyuSW1ILt2pHvcOkVwImbuDOPm/gaeoDVNarbPJhDY53qoaf+vrB
cGYxUAOCzY38cnvXVjQiy9oR/Ri8deoABegrfzZ0SdWGr2/m/BwnQ3asAg79jh0He3HSXNkWQfez
M09QSiRVRnRRz2IgpUeb/MZ3qX7OjgqS/Whn7pseMTZrnW0R2fxrDBfFrRGqVrZpamolYDPRDRFE
5YVJxRrYBOFTo0+clSFjvZuqwsGwllGrhix/MfzzXwEUc3jnNFDB5BQ4HeHoI/CWHcp8iKzbAin4
nKCy6BhII6XYLm2S7M2MSvvMIiNjjB3/AsQYuDsiR3mzZ8Rxn6i0wwmkZt1ZN/9zQiF8Y75vqZUU
Fyh0lGIy/ZD6MVJTmHbg45405qCGFelak/+q/TKQPPLELyEn56FJc8M2xfrnedwU87raODNi+Uod
kFVzBGBfCm4lRie9oSO1qnvAylL3xSQn2grI6ecEKEFizgj17wYATmiSzF0bt01LDkIYavHP+4ln
cyaO18Ofj/79mBStASAEneonDCz5U8eyKJo7A5xPnS01Yrsh+xyCkaqQ6NsNTBTZDuXLpy/16IF8
wFHO1hQBD+wipvPQKSW6cWdo3y2jdHUPzwC/6hPGBMXYvJNwudz7W39yDmxXcaBiF8MaubjCF7PF
/ndNHjpAo2xhxXLNMUKKlJ3cEAkQlxof5FZRJxb9KXau2VqnUuoi0ATDmq2nliyYmrg3lVHE8Rs4
ORehY6ycal1/3Pk9wXd7okWkpqLWVXJqiRamoIB20sWDl0ijB2IguvFP4r1o8bqJVu/aSLfKu3MT
nTud1V7fSpxoP7r4pGj/S8SW3S+ET2HSuFmbaDEKiWz+h+v+hS0GhWAbHCzvgZpvKTxAUW34faY6
oO90vXpC7bsZCirPfuHlBgkS0sFrrzF+bwFFoVxm1/buXeK477Cm/+KDCqZXeXbv18RDbaqE0Ja+
283wXAfevyvGgMiL2nPQm4dD1SbyuLAH7tLZS674KQG6kulSo8mXL5xapUwXI3AEX3fazNQOw9aw
IIg42ktNoF326lVqC/FL1fq1yMQdVRvOdZNmfEb9a+m6QQV2ea+m0ATRQXuCBfkFONiTG8nq1weZ
OfTXVlT9VkfdtsQbmGvnDF1fNX1A2sHIqgo4Io40qWmzY9K31YoHB3Lwm4ws8yp32vVtERi2sGkV
zZeWniM1ql42+aNTDQvhuVDU+RxJhu3h1WZHii1PNkj21RzYJWSlzQd7s/GEDu7vk6FZKQ7KwAxQ
WfjK+sGgdlhjAqp6sHmB0eWAbO0q06LceXjSbGOglfe1y92G1jtE3m1DVei/fa/2Dl4U13erdQbH
lkunzpRLh1CaV6ciSbB9kOUZ3qyxy7w0XxAQM1lwua1i4+QsK0KWW05Z8ktnGqwVta90wUfxeXVS
FF2F4NUGLziFRnVzEvK6dNTwTQpy9ayka1+TjgLt+pnMytlbCtaeSKMUhOqaFGL0Rj2C7xJO1NVi
+QD6hJtgPX+BaEl+Okk7gWpncbqaumjvK6HCU48+iQha+V48ikj+f+N+XX6G7sCasXcNIPI+Atj5
TcgzenIK1jiNhOm62n+Xu2TV6gA0wRI1LLA/g9gJxy+xwgvx01NV0bs1iv/iSeF3DvgUdB62hctt
/Dx4g/w+SwYwJ242DoyqCe3fGgxW0F4oMvfzp9Ba5zLZqBQwtWitNRL7vEkbC1KPJQASxbYmVNLT
WcRN919JuIDbZFjcgiwyUcNnbqEOOhv8joasmTlYkJiT9hA0jXgYrlcjsxI/c7orZzr6UAPIkrJ/
jnQ1zGr1stiKlPYUF4hosetoX0wS85uZ/w+TgHT7ajUQh4VwHxGJbtn4/MD0ZFEkFF6evt0v7mnU
wlQprXgPmEsgxIF9vq25uYSyLkY9S8Xu5UJRhB7bzE+W2O5+/XGzMfOyHRAq3Lyp/HAqryGeUQiy
UASwsQKzA7PdqqYnwizOM5+BVt1v7KvKRcdTPev3HtCNLILMesyL5MK0YFVcjg9eektZBsTp+Ao4
kiNGBtt/Yl6iguxx4LAd4YrmY/7b1sVQyP1xJQoVAuGXLJer9j1SScBbk2XUeONvIycXpyhbH5AE
uABWDxZlX9kwB0qdZ8Q2oISKKjuekMUpieG99QpVxeq9iUuqvlWm7R/Sxm4eK1hUCbZ+myEIY9Zb
SSWMHdmwVeosew4QPOSH9pLCekKHvHIZfPjye4SsQ9fJeYYtVUGCKWLiydStI3WNA+6b4b8q+UKj
CcPQoun/x2UPe4v5XI3dyTFwmQBUaCSUAxUvjoS7b6u51XSywaOC+rNfF9Cfl9lRr4vJp76w3/PH
m8gmVFD35c19XIp7KS2+Am2Y8Q7G0pbAsbLT+JzWFurkdijfNyDyHZAZhHCOzx0tY+p3jlX6hkes
NSu9Yzgu0LPDUWM4h5aOWuyVkSCiMHVqjIwYat4JapjLfXt8EYKK0YQ3RLJ2cQlbK68Rs9hXcswJ
cZtl/uScmH0w4ubIZ1RAPUr9+gxJQ2VwbixtW8AcNCJUWqi4raSfGUkmjFcSPq7oF6+ZYleFL71e
fQaKf4vipnhjVcSTS24cl3y/SWAImfAjqsvott/UCkhnCKM4l3uFhRYmIsTUdEneLiGcbm29TUnB
VM179/BQOV4sCt2VZebdzb19oEgj8gs/9MJb6ZVf/ClJZeDsDo24rdxsa/8xm1Rel1hihaQZ+y8L
i+iacD/o5IMq1pnLXPby9GoqnpE71FdAMGAjDZPIGCHK3XD79gdza24Qakozo54EFXXgqzaM1UbV
av58to7R5MUU/jSfzBVF93aW4V1/Yyip7jy4SicM7ALtjhaOXW8E0H0Fk5V/b1IT5p08Yb0MFWwM
vvHQ1UK+jyes5UNADltWOvmiJ89aBkt44VkYAp6ZT1hF59wedObCQfgg5QJqD9M/fJ3ktTBW366u
a3d9aJoPSr2AUbRU9SzDDdpnCP92msL/gGIEKZjd+BlRXl5982b95LrmPhKakM2O+xyDsUanusKD
NP9FKBtliyCiLO4cEo21seG72AD2jrfCsULqr47rkg1ps82VlbfWsGdmeWWaabhXN21RB0y7bHhP
/LKmZJAKTSxwrcsUQDGXF6o9R62FDX67dialiSsbMyQqJwp7ctXFI0KO9iZ5DnynKax1ndQPMbIA
1qZ9QduZ1FgdF7tSqe4PwhTfZjZ3rDkv2Jcp8WPx0KnbVcs/iGC9IkXASsRp6VcUHTlQaDvy7oWM
yJNpWtt5XCYoE5U9EUH6PSGGjkcE9F4D2iIqUKm8gOjbrK//RRbR+yj27mv7aeUE/pCOskq3Hhdj
k2AckDEnrEGWEAZUR4kU8GhsUMFJZZGK5gLWGpgZiVkmlnornU6D1BHvprBLPEZl3i0O+V9sRk3x
viTJqrgLxnLo/qajeL5ihK2RL70/pGm+0R0KxXB15sQKqvAs46Ce01SRA/MPzsP57pacCZD6YdZS
YGym1yaT9kDgHKOmG4P31OI9/aGs8FqXcf8RoMTadtraxmlUGK7L0e/GuppRWvrFFx9HmA3hLlII
8n+uKvu4cnrsNmxDwD469jms0Yd7m6EGK5xgOiNZ0zyHseYeURkZ5xaBMsEYBS3HE7JbTmpN/xVh
u0yqKJ/JoYQ5RPtHbXpMQv8LLJSoPN4sH5QCgFSJAjFXAFqKInh7syJcrWfjYumw5Fjww1VbuSmx
RkzoYUlWjf8XWy+WwGZyUovf3P7B3fCx56bsku/vKsLXl44GV/ZDrtlAFzU3IeDiIiYQa8JkBVqd
pLegL/NMPS3KffuSDBv7YvJ+bKRJ5LomDbiaFcmZSXxuBY6Ulqr8NL3TQERIEvu5oml5+ctRsbsl
Kg6zSriygZu4AXg3hTRBH4UqgtEa54w1VpM4G9h6dagrsGOdqUYH+VKnpkMmzEo+QJQyeaCt20mU
myevN+eW1YC2IDRXRl7iBs/vkc+md9nNpT+Zt4pxTJi33/sPMFJ9mHvwjCI3YdO0aXOnFRpqt0Mj
+DodaIsfZKoF/bu1v7fpbtFG0xQlaxiRb4VfyYJw4dm825ERpW0k8Eo2qDtZtvGTEkF3QYvOmLz+
NWwB0X2nMSgAfdcdZZuIxYf+rAS0CgaOjNzIPlT7gszeOGd3ZYgE/PSlDO0GIAs2KTvwhQXaFskx
1e39XwQceFhkVbc2pDTse90epRo2BvSTYV3+ClyG3vkA4atbsFMbjlYOd3Gt3DsFkiWEMagszlZk
fSPyzOL64WpE/YH93pA/lT5ICc0632kpjeK4wYYYYdKRXEjSSunLb6PTZTG2hozfW5AMGdaaADeR
chzTqX0Xz+BX5+aAx/xuLOQQm9hFdMWX6H/HdGQUxBauBFtwISzLr2xntjU4KATyrrrGYTyQon6J
7fTSQQv7/xTpklII2AeAo5Syv/I2FS5GFW/SJJdNe3A4+90DQnOC2qvP5iDcIYx5lGzvk0VGJnxx
C43DZbg60rpM0VQmklWQah5YOdAfUbGCO2p63iWmIuD5aVPA8c1iRoYLLVtNJgkifQr99ys+2Ki1
K5nEbdBjnDAZh67VsYkYiJ2ubrtmZ4p//joNARm8VuMmwewbXuesRmS2nB67CH7ckHRYCz9GLHZz
QM4jklNzRHd+Hoin75zgRx0wBhbmc2IIx+GQp3ulMxvTlbJO07sqmBdfz+SiM6d5jgHr7AQ9mZmy
US9RT/09+ZIPRaQG12nkZcf2xbkeitL8Ok//tTP0RKZl0s+50VtrLvg9DvbjEkE0uL6FKun7FwYF
KfW8BBe1AZo95RY03E7mPX/NWAiEYvaEmKCBTVxpqN9/ELn9XzJl2Ytv0BZMUWrKxEkDnTQIlgWz
P2u7vu8WLyLoe4JSff2rHPhxwEJbobgxrJII1grWdgHAtsK9USOe9gdrRx8mqQ7wUqSTQyg7Vimj
LOpvowPrHb+qp0Dv+iNSHRLIB6HzesuWJCh3molIoG1kBx8eWLGO+Z+Lny2PddUNhCiVBVcQGauG
jWSAEiJum5GGwNa+d9FFqoyD0/qpyV33IQogI1GCX+CqOUHWh1KagIflJyDLj+ywAyUszVBW9C1z
tECgP0nezDoKiSjnwSjXA/AsUGewGJCidSXTGs3fXUizylbVQS/CYIu4KrYi/AnksWFYItkFLKRV
OhOQvrgLVaNEBiHYIHFYmgeHg9HuBbVosPelxHIsj9Nxk7psNdYk05WjHj0mgM4Xmovp+fw0oT73
M5F0Qg4xzwyhsZktvUhTcPjU1pmI0jCh1p8/sT7EeI50TW89AOvK6n8IbpkzsezYKytRcnWu6hBZ
czmJ6RXZ3mbZiCKk6lSmFFoAUPY7uTTHiY9YPEngPy1PAF2vjGTzvjru57Js9bZeThVkLBDWRXlu
r72CD6uJiXxLQO9229FMgIDaIT86C8KKDQObAW7457JyLsICZOG2UbmJaz5u1tQosS2vEpnOgoYs
BhhDQOQmh5VZtzbJ2yPNDTj3xTqebegszFsSNnfT6ujlD3Yahttuh2J2Apgs1wuM8t2WfRJOjEkA
gfM9LkeE52u4O0b48dmw2+g/bI8G3Ax+5cqlCP55C1A914AI4KyZvCk8QplgJRNXs29ZYLH8hNDD
gWtwvKqFC/4Is7pWJfNGYVY0DQriDGrwWuwhrLLAlokPuZ9AU2a3ylnX9ZTdXWUywb5KUdbCq5Rm
qw8vVNoYYEBfqYY0SDD2AGGgT/peyU3K4HF1UYlnqrIIoHQ3A0wuC45AUFKfqxqz03DSpQggMIsI
1adqgdeZUIReufoH6JJY+7Y7rFDD8RAFkjpI1Fj5z050hkkRRRVeJgBmdG9O3Kc1ihYTaQXNVbhU
McxKF0n6CsyIrSj3Rj+o30yX4Fq2y256zHAHmG6nyEORHxIftXoNf1cLp29zaI4faQFQ5QHdsCYC
RFSc8AxADhKv0g7BujHPjbOpt8TXCe5tA5uMStKPpecDNp5AgEdHICKdpndgjg2TPWHUmDcVxwIJ
zNWkId/0vHLiVrcofKvufPh87dxYXBgJraY0G8SdMalQgMWxhKCiZs/OU+PLNIUvZAQupDKw/kXd
c91QMUi4QAb0eF0Rs3iAhVYrNbnpNgHnuQuZq6ZGMQTjM8QjJQ08QlWgsxDTeqlDQ6uyl6O568J3
Kv88zxm8zcEjF71PRROvTBCgmizPDb5jqJG3QSvEFjO4raUImuCd4YpOkjjGOf6F//ZqJU/Mtv3c
uPTLFSU6s9pPAP/OY/HWz1ByBjG0+gsIl1vC1prPr01xyJQJocpa7nScIvp+yj319NHMwHoTJ+v8
vrFgKBX+05fRfH7jrBAQ5DH5H33FTCf3YlQYhxeFmrH1d3PiUrkzCHoBS350lRYU/G9+eGLsJxv0
Nk8YI37/DvpPcrRgp+Tt35xxfsCYNHNOYxTAiIhJz7H8CfnjG8gzqzkhEtl8JcnkC1h0XifCIRJX
x/LM+1MbPs4kQdXin9SKc5HRW9JwGD2Fg4hbnxNzos/Nu/91j2GiH/YfTGxakT2N2jq+X9lIkDqA
SikqCqhO/ASs8o6poEid7EYwbAZin46hKvXGu1fENTRhe/hfa0IhhzKRHEKosX5mq1RDlSpfqadQ
aCbQs7ROsbleIE5ynbVWH+RkO3VTBQ+7tx6HMHmjZWSSfExf8tvYUpnIORCqUmHdwcZERg7uSVnE
4sojwr6knOYFRjfsfD3PyPj4f/uNJFlEQXbWPJn3MtKBeLENJkXNfLxpT5X41aXQeFwI72Hdgd9D
oMB75ihxCvSPh8Dxh4ofJtUyC557HZWMwpN0UcwTKLhw0UsV9lLNmuiYdovg0T59kcMzdQUrD2HI
3n/yM8HCn7z3NvPbRA4dOKVxIVKvhl8CTfeEmKgJfsv3BwTMjsRhcHMv3CI/kErP/h3cuPNll5ys
zWB8d5U3Fczl5WwdVhg7hcekAqSCWPqAl9CcfzMXHvvUzebF21D+kqsW1OJFfnmNNcQ7L6jLvM46
Z0GXHLIWKGve0FVU6ZJD7VJv01zVZyEm129CIxMVkInif+VQwot+OYOxCPMz7xPKy602qKP1nEHx
vEJ/ScxpC3p+q2jHFmo0dPa6JN1lNEwJ80bt9O8mmj8Nec8j6z38U/ih486YUU7pRqGSjldVJkTK
FuwvGjPRCs5HfHLT5+N/EdEVLBfI0SBbVJGMf2mR2SY0tg8nnRkEef7t1vbxr+5V7uzSkhak2zuF
UTl/6PPPIGIL7b28ieo6HYFWhLcCNUVYB5XkAP2+eobP5jRh53Awyp8peeNUYqZ4LAwbCl00x2ej
iYWSfWBatYF+bqBR0MnV2J4v9dm04nIaYk8ZfFkftIcOo8OqjSVpBJL8Kc22tcMhMjTT0zOp4ABU
RqAMaInURzThbraeyNMzZncWkgzR3UatsUfXLtqYyf08nIZqkwNn9JGWO+WZ4TRvW04WoTPsfdw2
IpBOH+dctQn3t9pdeAyln2LECuZlamTHZjGsgHmUZowgAFTjIAn5qQbb5f8bjk57+ZQZTWLw64tV
FOhVZMxVseByLs+NEihet2tVk/RA9CkvP7nqO4vVRxqOwBIa7pBjOhHvDlttYmqG7oRng48ZLQGp
fWmNfQ1OES7h0mExUoZAHUlIEVyPVTSDQTSX2X93Zov58LhT5DEZB03lEMjeAuQny9XLZ17AaQOj
v2C43hDlKvTYyEdU0v6e8ZeG72f9odL9mxf0N3Gs1q/Pa4p/adEMJOKj8wwie31c0wz714EbSutz
5VsoBeAUBBM/jgwl+ClVnWoNJuMLLUeYlgMygVQ4eGuXK3+vFQLmIwj3EuwaQPQ0E9P8xnIwS3Qx
1/Ri9i8PeRex9s9MmBl/FTyP6uY2ws9q4Br4JRjUjPhJI7UKVrALGesT02sRHSKHLWCI191DYUq1
qttZN0E78Ljx9UA3dgpCarzBWPNFSPYFtAhlE6oqcRm++U2g2jeoAYG1ztLHrvtxaaHf/tB+DG9U
r8JgEjEVdjjodkpI5/Gq856mBqOC7+U+zSTS1B9eCtqS3rVj/5vwfy0dwSnw1g5tYcx0hNJ671Oq
QNYFkF5BfQ2W9yY3fBhic3SvRIE7YtCE2/xq3zywKQLQtto0IctYSAMcMEY+Yinxamckc7acWsCc
3xvZor2D2TEEYIy158mAPQg8p69B6D+xICYeV+62XsbYlcO/5anhIBmTDgX254DpPUBuxAmcb4El
X/xL/FoumLH+fx1/fMamQDxloqy+Xu5G2Q/xPCWBSghT7orIwKI3THgzw0SYgURDNexIu9CO33UK
XCtFiMqYwks7l4cMogp/a+TfEt78F8eJpOoXLajcr3JTdUBwGFCLiUJ58in7PBJl9oOcZJIl3dYY
5Z+/cb52SmVTRVEWLsxJ92a9afUfAjMAo9m1KZsC37wq32x/ZePVcec9nP9S839jnAi05fL7qJkv
nSWAdWI+WM+AZ5vr/h/QgNgI8sBEansJGJEAewrV13Ui5tp7dyoiOOnuefInSET2Ao175qwfFbhP
qRjDWHEWO1Ekull3cd5csEUiJsW2+tvDCyYUK5So7ias6xzMmF98c+yT5ZjZt7u3xCklmV8/JU7p
UNifYE6BTzBtjSbk5rcI/6X+6laGD+uXDs3SEJdgmyF3RYIHF8X4TISatlQ7QFU5oldqxBQ0qgXP
+0vnlQ0Y07iDtYh6ue3nBSXnzkvo+2c2IQL6AOoNaMLbRS+pNnmEYkel1i9I1SanGMvnwYif5f52
wVs8OSPs0SvRBAuFgdMp6nReA8LFuUMaLNf2kowreh5dOBKmlaDqGPpClujTFHD2dWUffsMNypga
D6wBchn6SDg5L3z6GBPtBbRU97JodmYYRnU9/KHlBQIumkh4IHzhvzi6Q9QDcCxyEx2v7/URHKd/
X/+7N7qD/CvwbqYE5eF/vTjmz4cfJgQcg6OL9X0Z5xlAF15vkaER//HLIxx9uben5ZwZ0npqvblk
yOWbxwveuQwOJod7eutkINgaAft6pLRuAJyeQXvKXKKBky7UU+mqvBMQRI5FGu8niy/wFyR/me28
nNZwlPebIrvxJPwAVE1vw9CVPVjX1+3DPwIAWio8WsI6E72zjQ/hK13miWXYb5lbx5scXTyqdmZM
6gEg6pxBblBC0qmXNKXpxF9hIKjCJaDj4AXuzHJpj/qWFofOuZhvi5RdwgAPIBfC6yjclaKkcNyS
exfJ/qKQ1Ux37sCrpOBwB6ga0+kyQrL8zRgSa26O71J3ruXPIr1+dQVsqgsLE3CgB8gGl0RRShxK
N8A/ECplUhV2FBWgtzDYCOQEKrZC8NU3tZeQA4LHHgPBcgdMgeU9i9UFA/RYDl/8nTmLV1ykzXfw
XH1gO9EvYbeSjbJ/tP0wbTdZZZfskXQWe3e9yoPQsxSifym0ZxnafpA+uzfrbBu28TJ5yxTkLxGB
ViAgLgB7EZ9FVh5NF1s019dThw5qyNPHF27jsW6k5kZi6LxmnhkRAx/KZnlCk2rqwhopS7wtln1Q
VPlcYuKmmWT6dYk/+usgWoGpoFxMoIuONgYDy+u6trW4OYDzLyFJJC2e77D5aLDefppzFISfUd9G
FhABKQWF6H69DCZUHl5ZgDfwls/wJjkJjXUvQ5nsK22euN38tkSp/wV6OfaKNoxRPlSAEAPeDUPo
fE5H9hOg1GVCkDaAzrOPqoWeWJ0uIEvwvLTtSxSpv4CCEl1T71cJ/C064INDpfoD8dkhu4NXj7Lp
b2KxbNm8GEhuN4uQBRpB7+RW3WkjK0meyX1ijcrRm2h67/YYlksmjze40c0LbN8B8zcRIB/8/Pv/
LLhtNNSywNeXjb/MkGuKiaQkwCsYcutImJqQ6cA8XHzg5gOw9D65AscOIxdcRtEP/vAese2CATV/
MkEtLpRs8BdaX0PgnePL6a7H3+1XBrCbcutNKa0F/gxZ3fpW6B47Erevt3ajfyQaEcol0YpfvvNq
K6/bWDfnQjZXE9+Pr33DBWUGO0YWLe1nIGAce/gPH6VoQgBOQUr0SxL3gjVemgd3PxG7Ao10MF6v
3Xp79wTCyYKdfMGUgofTRQjThLUTX1uSUXqP4m87Wava74Oj+hvWDmoQbGjcdfhcoT3Q6tiJ2Tfs
H2bmRYNrOAyyS9NdwjtS/ohtmwmmq//+4iXMdwV85WCOy3fhXJLbconlKrufmmwBlv0866n0SRkP
yTBsiDY7KqGkAD+Cs/zFF01UIPRDI9hNuZZOTXONjYxP9MVl0p/mGl+KHf/GMyphQ49ralY7slPy
oofVFWJvmGRei9pz9YylH5YQFoMZpE9Y18+b6kHfWt0tSGTn/Kf/Xi8SzlVICQpguYrwpw1qjbHZ
4wPJpEVlqlhKi9NBt/0I64Ebpz6kZLv/5Z37DBGWgx8vEof5OMDqXQZBoVwTq7KIX4XBHgv7FkKY
m6N/rRIvTIPk75CJ8izDsSTRNDXS+23GaYkUoj7fwqXd8MadUFRkhtADR9+21zueHtbpcRvQ/cpU
NXMW0HO3VKCDibEHcb8R8CpbULaNkxENIB1o/4f4Zck/pG02r/ecek01wSlBleLdDScmx5Or5WOk
aJ5g03oSQD/mRg4X4ViC4h+MEDC4V9k67M/LbxvtzWN+mhVEYpv3yWmzr5bGJG4CNXPm5p4xteNq
tyMt+d42GpjG6b7UoG5758QwbLi4hCmGQCVoVP6sASsRN2tRoTyPwnsb5Ch5gT9gC2lItsREgVKz
dfJzxKTY1gBm0VcrI0db9ikTLVLu8KeZ/BQgLub2HQayMEFrDgJsP0z8S9KEINmim+Pi0BnxK06L
/aci7dAlePjDdfon7xRNyOOPYluRRdXakdmp9yEQ7Ug4y7qUw9lFRno8opVpFBgSmh13UiBR5bIk
fKqGN3zQ6v9bbRjsfxnIzd32t9C8hIoAfu4Xy/x7pfJuWBxOdsM7G2Zf74oMsaE0yj6Rp+mQEIJp
3gbVniH6uyHwg1RkfeizC87kcvXJoQsKKUgRorOrZ4EG/SA/tat5Ii55OIXE6hapxFJCE4a+jL91
9eA2lI4qEWkjgD7CbPuozXxuftK6zQnwX8mI+eRGG/FJZexbEo/tk8+FWddDe3l9mPp3yQQwuQeF
zCXbCBGd0Mx4KONGWGxONCmX6O+iM2tFAil6vIb8CJ2DCIgTeWpdQbhWMW3roVloxRV+sU2s2Ahm
pQWqi1k/noH6m/XMxNfjfjaiuScJ7TzPz6QWYH7mNfrclaYN/B1JDoXD14vq9lGkbvQRs1ZVxNhN
+V9UrfmW72lcS8XfifR+VVJmrHZB3KdMaEZbCHSJ8zzu0NKKY7ETtGmbWfI5gYR+749TEogcXXZu
RsyZXmslLW6mHPsoGGVpKuVehDjurbl/S6TbPar1MLWZkIZcmjg/ZWXfO697wWJnNdnIw9JtDd05
dmXTrL1vJVB4sz9I+QXBMyYP+m/k5B0fArbb7r2oq9wi+9lnKhPZgAB7JAygJ10jzeaCERccszUl
kIw2BhpR34GjsnBFIKevkZLiQ5ZzjdTJ1I0HeT3HBfBjYIKhWTToZvpsMilWol57DNQDVRjRFZJs
JIHeUTBSoUDHJxLo7WToJ+nY1bOl0G/Z9Dle+7goDR/Xdawhur25+9xPX0BCL5eUWLRbP4wGSG39
VnqYp0USoJrphDELKR7E+LcuWWh+qOgWwtv9C+nw9L6ZHe5+t88r8ESm1Q6Z4nNt1DxURXGvpgMP
Eg1nzP8vlEbDN/YrfW3ao5rfEztc+DaThas2pigq+Wer8OuXdsVTegOSqpxjybe17aqw0ZWNHJSQ
4DOXSuFC3qG72AjaQ4TyqkCBOjA9TGo1YlbtbqA9TeO+pTOa09hM0YOdglLlK0bC2S3jI9Bhkn5q
a4majDXRJ+eprpefUR/2tQf6v23BzMcXgtuKfURD7pYgCMXmPVhUPgpWsi9Z2mgkeiXeUYv/KSdV
3+H9e/V9rEFjgEEm5YqvdjY7psjY2njeGH5VvdiAlv1QDa3rLXgi5vWfJr/C96HiIa74q+PKAXjl
zI/YLHc2Zy7nDbno6o6ezFbPKMrf1btZD5oVq6oFzv+m6y7SjhArprML2FqEO7DP5CjJRAErw8cP
Wnt1pN0l2y838lwl8G9q3KK+Xp9HTb1j9M02lkmN/Kn9p1Q2gp7SHfHOBgzPwlKnMdnnOaDiJw+W
wxhX0cTOE5YCj3scfuBf8NUKz7AB+AO924155jt3S1MlzpIVmMSzWAov7EEAvoZUnAOu77/5E2iy
27xYfnq3oGA1dh6wY2Gy1UIoK4fh4U9B8v74pnldFQS3lZzecYzZDiWBBbw9gBSeaxquTqo6j4CT
baFe40TrN2IHCy7nByH4xPnzYOKCgFvYkFJZug2tlBvA6Q5sRqcbzQWZj/Yt7DqhPqeIfjU3cEAK
vp3hmsrzGEJeF4wjuh2Irg6HUXNyXH7Due0Q0nUPSsV+SwKe1SE8TRQuf1dBtgehs101KGBv257Z
oubuReT9e0y9xmvxYs+uQiDXc56wYLHvxpWJo08/AK4ML1hZSLD3pSH38HTuxW9+7MJEqbqzTuCh
PcQl3bh6IMgDLV0KV5TLXN3LpZyZ4nk2r13gXHB23TxyARxiaObTE2kTchItSDsr6qELh460VvM5
iyCC6IGfhhVtcEAKYNF20ciN+0bwrZBvsroE+oWNyji74BWzS+hUOT+sLnbo+2A6HbwykQrN0Vav
WeuJTfGPfde1YYqOJYr8MscyC3D4chRkmxQuCU62CDl7+tShIEH1obEP2nDksvP2AfFlBgQma0/G
wLB3vsyVW7RQOcVJbeRDcGrHV57a8oBgpXfuSb64J08Ir84JOFjo5JBC61oQ7Pue58vo1IpmLIMr
qgE+QF8y/vRp1bfqUIaAo22Fa9/S8KCtkFlDKTnH+mKC2nybBreEWRfvZWcQAt7aywlO+FfWYF36
l4JDrCcVcLVLn8HEqvFUD8r8CotGb+Oyz3n3og8kpW+PunKdry8rDde5TiY5JVXSgOMpShwdi0U0
27FXKlDna4lTdF91iNMhHO/y7SnCT6upxvyv1s4IApm2K2vi3rP6PY7nDoQ+LiTzhUBgmCWr1uyY
N0AkIHMjmI/7sFEnOWSEsKTgsEiVmG1CnNxT3WQXfZczLTveJbeGIozhNZKB0mVaxr7zY4DW3+x0
AtNuJ1ej/8S0u99x7J6aTDsaZGMUivZrA0vAyh1MiMr4Lsi6U4eb09ri1NQFvTLPnA8HWL8JWqCN
EuuZ+j0mkz+rsAIl/OShZrF/I7FLHswF58mkxBYMjTqoWt96DHfinAQXEdqtJymu7v121+3FxUbz
F2v7KTeNGUFIkW5HtoB7tHyDUIxriBuy9e0VwKaUr137e4nb7w8Tq6BjnwE9VcQVouiQVuMjPkMa
gF5alPZjmSRvph+kqLeT0soYCrGIdNVCmP0koZDTfty25IRzVWcYzc2huTo5VNBiIAQFxNQ8AYWi
9KXi+Wccvh/oD0ByMBQ2oBvYc7dAOt5sYHBMN2knV+v4XgLvx90fMWC0EppWWyqRViRlyX3XwHU8
zeBO4HUZQ9E3ekSXo+3JqgoOYUVqh49ZRNQW7p1o9iA+xbtvIbG0AGZbim2ak+2d5aWqnhCvaqCj
MnPDWxHwDwg4hoQiAMt73iYUgDcSRL5HR8hlLBbpYM3VFrduL2HcDij5D88MBoXaMZwho1JN4vnt
YOdAyw0rxxtu9trLKpQQJrJ/v8hqQX+FkvyAuzOsJtfizrqYIVnS6TyeDFgE8OvOVRoJztruO7wp
X2KDDVHRCYuFP9o2LX5TTQX2Sxc1Fprrckspq2J+dWz2m0u6Z9BguEfAVfY2FTTXiVYrXU/Bl3f/
cN61AgGQVQNFVVuQS81bsSSCamFu6CZWAMcTn3M3mbZvXC9ltGlteAbKyqGVp0WGnTzzEpqZbEh4
FTF6JaQS4jhLsicbXS5Hk8mkOamMPjEKG0kibe4iUqGK27JdminVrDBWas1MNlxltuLuiEFG52wT
c6FCdNqgqH500TOO1Jal7ZVslVXoHSCW3vKEkV80A/5QBQR6h48sxAn+Li3mCJY8tphRj+1a4lDB
RXaJ/LQw8++ikx3YDgIrhNKVBiVnyKSmL2Utpu+9R6Ee2Poyv0RdAaP+hPh1Y7a+as9fxAROcMPs
rdhB+OTsq2ckDv1Rwad5L34JYMtEErUGxWJ2IsUSbA9hblQbvOGhYjRfiQvjKlgRtCbukCr3A0sh
Xd4Y8UlNrkdv6H+ehanRLx3F7AZK+7kNQF4I2OW3dbiWL8OUUnM84p1kXyyOqgD2WSuJ7FkxQZky
dsXBHAENO/XPIbxVQwjKyP+CD8S/0tK4RRSSSLwD2fyKykgTRlQZh2poqF2nO6MVX0g9H9+rOYtU
/4E6RvZrfmqlWD75GkIXimCddAyQwNcQ+GDGiiMUtFYx1v9Rf5D6amV/hc8g9LC6oQN8X7gZQjwS
glbg64WelTa84tQHDvZrV6F+t1847uNoIevTAW9TAO8fq3Ng6rFSWetKloHFhL2iXoEkcKXW+/1x
bVGOu7pqOpXTYXhV+3L99aqDgZQM7kJl9VkjLfvjJzzbZXIKEp+Gv3NNA+GYejgWQQ82nbbjNMGs
kh5JbIgokyrJZqH4PON7Yt5+f2PN30X2ywNsBkOgYPLRuGiG+mGROVI1ywBvYm8klBoQKpCbnstm
bWYmaocEjS/j0WTKT4Gd59FXY0/xqxxLQSVjA4GJEgF2eDh4pOudQmcPZMyvqgjXtnbF8CYCoIYx
7MYDt972MBfHufaUrOH3LmQ9Vc4xAeRXLZ2uQzY7Or3fkjcPkWQcQMJ8fzk6LBjCK93e4YFvbrvV
VqUwwG+HmdpQfMTyuNOgRjT/nEGxARr6/a89ZeJKzuAaxTsxVToMvcHzaKQh8EdnpSsyr/ZlZ9Zt
GpXd4aGCoFPvfbRwEcl/L6diEQl3Tg4sVcekwaqb7nsNlmRtD1rBQarTM+8SJP4CKO5T75n0kAVF
c457nx9WBRkl7HlwUaMiqYTodOyqOP/k7no4Q7XmYLdzSTXmdSD2xpmarztV4cL1sV84FabvM3t3
01XWOVAkrIALERgSC436NRvWwh+YnXn5HYlJJ6BstXa0/KBnyxzyXdmeRx+PQL3MhEtTkYG9NZWd
qEijgGnS0jg0bflw1/Fj6i+2tX1RUwLuHxBkviMn+sNSLWiUdd7Iljs8iouMWjM69zn+15n+BTxL
z51YZKcVEy4rco4o/fokMyBNl7f/3SEd3dvibGzpP7B4oG2KCs0DiDy1ON41fawWDZ07+Di/6OwK
VrqzFAs3oyPesVBoZHimEEdWhmYTNUxCxl0zZ/UMsLNoXNNFxTOq2QG0uih40Y40pMWhdNCYSt0C
4Zd8zqyu2GNAGRERLivyBra0uzGyAGTz3lrZ8Xq6q0sKt89l/C1O7iFqhtEZe5P5tdv9nt5SVGPb
lgzumUVtyhMQFXAdTXddWYkMGBzGzwPHlh5r/j1MIlj9YbaBrjaRqkQlsmlf7WdrE7PciKFMhGNq
DzGXTDD857wj8Kngtn2D+CZ1nZxZx3EPHf17D3orAzZHW/xqyptcmIPAIMzClLwSjNUxy+jhHi1n
UXaNdilWCQTrI8qLDw0+UNsUP8ejUzffrVVH+CxFYvbjVDc69wzhD17zNC5QMmnrp07Vnig+Xixl
jSFeekF9HjhJbxPVp46cPS8FkaEA4oq9JWYKPp797A/b7qyGxAnQwOSeFyOlE3YvJCURzVrONC5b
w05QJpHlnn5amsClrusptDQHp2egpaNbjEc8WzcZ21mBYATIxM4kOUDYRVqO7zskUxsxKH6bhYeq
7CzbOUBdLnFXJahWDiL5esPZErhjLEyEdIJffbMY+K6o07yvEXGyF3ZuQd+koSPLdHQDQakiPZvK
jiaQrX9RmC0bw7Rg17RVOMHy1jPMF/tk5x+ITLB+dKkWHEcrt593/M8A5+adWlHeq+2RkedZpDVr
CzPhMXzO4jY6P+o1Krs0H5mt6kIUhf6P8fup63EW0CCq19ymJ0VBqy45sI8HEMhLALHVGE2ZENq9
HSigm4oJ/4Onz7eFdVcmRSMPI220ucTDIQ999lUPm5yBejg4UTNHWKsj3ud67jT6iwWjv+YTI87E
me4fHOSvmaQKGvNj+x79+w18Zd6zHbF8IbJYPI0hsYTNCUDDhd56JVXFH+0aN/ywN1q+VljNwncH
FxBMU4ZFs/GpwrNMF2r0o/OD2aTrZRoiQNUs9oi6LLBfC5rRCKPZFV4Bc5DaegNva5S4nNoyR3aw
evdxhxBSNot6KEoszStsRMK8s4W19aPXgKPucd7sejcyp46P1AF3bRwUJq0HNKFTbXAM5lHi9hOC
+mkXD6oxy6yTOBXuiPjIjNqm2GTkTCj9p/5EZqm0OhilJeVYygYSCp71Z9xYhy4kE6vruUStkx8J
eZQZm7YXuvpVemeZSEgvSYeIma9d+LN47k45z5k045xw9047edFABMiWzANV3rSbH2pT5D8PlNUJ
BGBpwcMIRliDZfXJBV+48bUBJXYjBJtV8FNYwHLeZuRcGL9fBaJyULzjAMa9R4Ud/3M67Fwu1eWE
dQhFXpSNJzKp935iUuX9u2qRPDxpywl684O5xs7Dpan5w5FQSg/QuIB6X9OooYk4R1W3hI50sGvO
hehx70EcnYtZf7D8kz3sN8zDrxHSbZqBRLibVjV42bZUcrOEgkokyHXdHFk2Ckcifpw+uXTvivZ1
MaXiTN668Wd9lJylS4jF3tjkuWps0R/S66FzuRdgWm3NUju3UIhpp30VdZEoXrtKFurJYTM0X8lW
tdyJVJCR6VE98BA61U9D8hxepI1+Y3Ha6DrHlCj+P8F3fKIBivLLfQey5gHJBXp+Y8gk5ZU3dzEs
gluHfbSbzI6uaA7fmema555wdGZXxWzd0zwq/xoODCtN+aOWaiQmpX4GdpLJmgL2AmlWU+JacTRq
OPxYuBTX3MZHUgLALOphuHlkgFQ6YUd0qSbc+NqRdf6GcYrqNUCpGOxDoUsOtXruLVtHFc+qnXOp
k8bZpvsprrRbTTl00S1T8YwkCo2/c+6MkoyvwCUD/eA6GtpQF1N/tldE19PftQt+3XaDxyn1eV8h
TP5edQwlR9EehKzXUp1qknsLEuvw668fDxH3tUSAfqMrs7Ck0+8vfOxqZNBv7we/Jy6Un2py3GwU
f/QVMH30rhTW7C6qYV7OL/dgM2TxW81j7BNFYDpDrTJyrK4LBeJykjG1HwwQY1Dv7o07eIKI3O5P
6wGHKxINEdO7YRAUuOuf3JnGRUWxM+BrS2K1acWx9IOt2xpaDz2PWn7GQ2vHtY/n4lcpa21Ze+ZZ
yDbVYvvXyYspnYx2lObxCYzVkS2TABhA76glKwlSbWE33zdbSDIKI8/OgWRdb3bTh9CFxdREin1p
HITHEQRMtlgUQDZrssnbz6l0kD9VoGBjzUdnLQ/U8Yf73p/8QcR9gAj1G9zBIgMuLmqvSk0yK1Bq
G8NVsFP0xgwCuxixJC5mZgyGGY9FEbyMrXfHzTKaMvYj7kbu121cdKnLlKlrPCw/x7TX6gx79Tmi
a3IyzOdechR1LJsECxAU8l95uA+scujw0gjELKqBfi47J0LgYJMnJki7VaDM4UKMDPuxdRUT11AA
wZXvwkL6Z4g3CTyPeA+uLEPaZzBiFD/Ei7UKxL5kbcSMJ2ojEUm22QoPSzoO86k0PKteAKJP1pkn
OkxzvOkoH41gfFnbrOvTjeQgEVfZgUk9Te1xyUQnJF51XTFc+q5F4eCr1JtPQxURhaxaRr3+Mz9a
oGNdzFyf64mrOuTz7PcSGilhzYfC4spOIHQy+/4Sc6uEsbCs9WcstjHikcVyELDmDGrTENhJLvu1
z1WyVWKhA2OKKgjCuW93FG4r+3fz5uNb4TuuMIDnxo+9WLGYRG0fD3EkPPTj32rZ3YxOsl2YHwTF
Tz/USnNg77AMmRkncen4bx4G59BAgTziLBA5jloIRyBtbGhuAFquFUnbJOyuyxCj+j7FJgaFxqmY
AtRyKWxFb7lCCITTM8rxQj50/D3QfIw2WEUqKOkIGCBYSCzLGragl4pwpAzj9ESx84vOjKBGotkt
BUtzK/5VAf/fL+a9OrrRlSkVQTxu+29aFVeceyQPQAAyf9sMF2JWBRuqcsB+3UPPjdkhVfGgqRw2
IyOxtTn20J3HDJlg4ZdUReJRKs9LNFeFNg37AIZARRZTD5Y1oPr6Au5tDtDmFnK6fLpEND3TS8MX
BVk5HUsKedgrZ5h/SLkUbUyJyvV7FNxG4g+Raq5zH6/yYsYxaOCKE6dffCmyzxmkpRmtAFK4WHEJ
cxIa28BvmNzRycvD9+Skt81+fgDE6IsATPsJ3acgmx5//4xx5mnQnufg5/DlhqyY/c7oZR8xzoup
o3cr0FGwwApZ7QJ4pAo9EGAJTtCJ2eyajUHmTu0p7XRij+QN6KgXmkEkU9vvy4oL1GVLxclo14Gn
RNl1pqKGAgiROgeraaRFfr9oDxS7OQwPU6/g46Gc+rjEnuNmLppMBIeJv7R25bAlgIYVeDSejvdW
BKXjw/IE1quhU/1rOpBB3bVVIt3IqxMrcf0+RJ+5HkLWIB9pWWHUgkgkgiVlwdAfHPGV/wggepAQ
fcorTT/Sy8SrEz6jK4vxq+26zsuB4NjtziTyEwGVqzUUBF3nIZ0QKeQA9wOleXoB0COfYeUqmOcT
mSpCeZcKI2uxd2jfKOcbrQxD+24IyVWLgiGFJqQlnNA2pVSMZbjW4zLtiR8ndfgPuO+pGgy+7OR7
/MEcw9cAXWxRGKx+C0o/B8Aa2Gm7HzGdQGnyK+PaCpl3L7VgVXcBlzbwszR33qpJpev+CyLK6RIT
eY93sHXwrYF1FeW1OGzdK+tH6XvRO8OcBkBMvRrkTu9ZTUXfKaPNhMwV8sv2a7LIKcEMdCOIL13h
DRpefQu3q7U8wyH1sTPTNOhIN49YNR9Oz7y1EHikZb2KTKvEUhWhuNJGXFbsjqJZr9jxnlLkVWAs
AvNq5zlAHboai6oYsYJdAeKTCK4NOGjeUSF1qSGYhSAX9P25sMIdAyRmWCzT5LmrxXP8itcHvGfM
0bC2cyIXKLDLhPG94zGU2li5DBRUg08jXsbDgDZkwBetcQLw/y4aTahLySkibO77O77XB/9QUUDD
/MGlLiOCbTmdvuUnWiWCX3xG8QJ2Rhs1UFHrI66MXXA1G+DTLS3PRNleJjzmimKbcbnRon6kBKuW
tSBeCDqCdYvo7x2swbt+9RGiSbhVzKD0djZTP3z1wtjtsMpZ3NbAAnnIBHL5DtRMK3yIbXsZZ1G7
jOI95WGPUtRheas41jjDAp7bxa55mrWyWyDRMJl+cPnf0LF2ZccacyF+SRLLwgAAKpCWoCGRmqc9
+Vo61JM191gQ8uezGG58gDRDuIyZ2V7rvwnkjb108hcznyYSgdxoa2fkmF01nlVetvzOztdMt0iS
U6Ue/wyoPaoYQNnINp3HnyL0me7s84qfPuLTl9WISvndy+i3MQk7uxHufmUi7kyTxM3vSFGEQjWA
4fJi7I8GQZH8rbcoVI+/c2TtIGzL78Je38PVIt2sOZ0/lizFPaAqm4+v7YlcVhBHO+w6o5GxY12Z
wDaT+ZCST7KAogn8QMvbhmc7fHQQikZlCgMskM1m1uGwDF1YLbnn4Vu5/3mbwNqrrYVDpO2EV7yd
cjdE0oEHwOk756+a8ZWo1dRkVGckV0pBhQQjtlG8wTfKIx32CuuBw7p+GFdjfg1DeR8Nq9jbBfm6
nvE7qwhG+VBeRUSC5z78+srIJcgyJpCr7PQ5Etm4Efe/SgXTpi+lz4onjyxLdDeZ36E09BWp+vmD
j86zDOw9DK/7ztiNJLJ2vCWS5VMwfyNOPn+K0recsiP7SVIOjo4pbFBKIiBmzPGmc83GWjxy3/sT
E8NHD+W+T7fz0UHBea6YtPkMQc7cOkyogdaxA6RLc2e2ZCvhfWdSiJGbv+OArJtxd2AKK3fWjDrU
H5Rs+rDPf55fY3/8qtpPS7a7UjB49nr0eHaKTZ8HHzqIcn25kpxK4kEGtlmY2ZHWYeIr1d85nyxx
EO7HhaJUCQaH+o0tTuT4lgSSI5UFehn+G0TNzy+q5Q0gH9Nk4UO3XjZPCVMeVzhFYmujzE1jS3KA
4id6FlHBCBIjvXrjB8CM9VANfuKQmdifkyBQCrMwdn5qBxsPkDvCu3qV9MJt0CqnxkLD9f6VWh+0
ND5vuTVoqYz1DT/B5uJY9RvwZqo1Ol7eGnprg0S4H0W02WYejPml7tuHNDLGTHhiRWmFg+Ae7rB/
cjgzOuwPhcyl19YcLEfb+13oGIO23HJyBE70zRGiUCh2FqDBvVTvID9ao6W+9+RB1adLw6w9hbQE
9ye8IlwFcCnucD7gi9idZcBgS3CenfDLmEK/q/pQy2pboO62Wy6AFP7BjSc3qVGBSnrnGZ/isepp
HPz3cCEtnpCOVF+q5RpmgDciuGEvTY1qCmimLjBmJ9Q31PLj3nEwVw/Z6xNoJj2Ju5G4JK4XUwlS
ex4YGL7cJaHCXhu4L+eavYPkUDjNRJLm9nK4wQO9WwEn8+/rlDonjARjJFyAP9xh3dZJxB3ZypR3
5g26TGVUHEoRbkMEaJDF46lT8eDdB0FPK23W+J8Zyt/fFxp0SKqW6enNiac4wJJ5YswNoQI2UPYv
dotkAHF0GRIQnyW4tWanYFgz4fC0I7vAlBx197pjhzw2DnZ73VKRZit98C+i7qfLRRJg4SDoYnbJ
4kV3nkup/NqMMhzk4qQjB/9zAmsF3luYiYi5wZc4M8GUvL+EUxWfMkFEh5AhJ8Z9W75v09R0UgAM
MVDJEfLs3sIufrynaA8vNe2EVy201t84kneDJUL76+Tzlbt1Lhk3XzYwyLxyHYDzjryjq7QGPKME
9XXQBCEvzm6puy9X/LQN3NtCJbb50PyAhYBSYta3N+Wiz0eOM0d9S5kPUK+5W4d+I9kyqFTUxdBQ
tATKu7mTtvsyrXGIvrj7R6TasriQGhjrsUVBjL1kMIx+KLtkBwfaOeQ4olCs2qagmWef9bxO0mhQ
7jl9EKoeolccHw5+EP9gogxj44w8NiliLeocHcsmiLJblnKNaO7z56LdjWG57k26dl5XTHpg70p6
c7GY8zTIPyTXTm62tZNTahbM5sOzO8cY/MxsL9ReleFcJd6n8ut5beJgx0ljcA/fC2yQP+JP41ll
n2zhgBF1yLD098XC0O+6GtfZO4ADBi10cpToFXceN72+crmaJ3bZ+1juPbEeT7KR3JahLxKOXJmR
utXhKWr0xUI6Wa031pJx3+9gHhyC5JGJ9nNCOw4ABsyqvOPd/8ScxJZ5kjiPJqi51c+apgVTRP9M
1eHBDRPhtY0Ifa+nVOVSD4PWS9QgKoKmHOTGhoJeU5Ec1feWpfu31tMnnnxyfpBrCCl8nhMPho8X
OjoXF2/U1ilW8AWHcc91ZPOcSTIficFsMyBnHu2+coQfoqpi07+uJvvQtTaXpL6Pcc0kvvCuMXGC
pL4ZvS1QSn4FWa9NxPBzLucscs7D4UqlWbZQn4jzYO5WPpf9HdakHTunsaU+CqPz4SmveAptNZiZ
AJNvg8CrgFJ/gOsDKl1M8E7Bt28GlcGJhzWeKlJhwdYp6qDzQ1Y+pcJDlqgOc1PiXhHFiHS4+RbJ
0KFlA06Kf6T68It3M3gU3vQERLxNUJ88m8JtXthahhItiXv4Xy4op41w8C30KDB8okDv1r3MHfO2
E5WTcVbC11UOnsq4TCYC4aPqMcjRszkRD8wYnVpEapBoCIY9VOkmou9HjLCtL2h7Yut2jmjpj4E+
6BSjbP0EZDMi/1rKFa6PpMEsrp5P9n7pWAQaNClXXtZLsMH0814jrbaJze+aqEjTfIPv3dhytJ8q
dPuq2TJcNgNhI2+KlTUYZnhEW4WiRuXm7QsxgDkKO676F7+mrskjLfcQ42YilPnbRgFQ/cKB42ZM
N1/94vTDXLmNIN5/J/cwK6g36PiSYpGWaN7w8FV4rBhiVl4wKhG5PW1vS1+yYnbQ5KGXMGJItSLx
8NlngRHlHINm5qQw4EPa234dNeHxgRVw6Q8XYp9NjVnm1fxA/HDOBQWcrKZspJhohKHq964yIOeR
v1vVU4qftiFsQVqV2s5x4RE12i9bzmi1x65pS+63tnohd/EXOomcbwXLlvZ9dLvc72Im3shnL081
TzAMe91Msw6FEfvKRcpyvgs6EQsldTM2DAITLyKFebhltKxY0/QDik7id7y/2emUSYaoDs0WwkIu
NO8VpMOC5UKgU6/JayNZ3oFzR0UaFprcrUHLzu/vcgezhbLDkabOgH5dRR5Ht1V3wUi49IYW6m1l
WHQL9H+jpip0KKFmovZueaPWbpx8x7BpmJh6dZz7BfjD9CPE5OUfBY3Cz3VuMR4V5L8aC8LLTEGt
bvbOOHwARubV7cyd+HjzhpBIhEHv990np2gMVJKBQmqMcxnDO/7Z1US9PCODud5HY39/Lsx3KYNA
lRQuc0bEQoVY1uKBfAyjrJKenCjZY/CD4d0dL9tYsqhEJ9kqsKQ3iVmBTq89UPRhYfPQDbfQMVsl
lrAEVLCDjFkI+DG8Lf5mbtYHIUYhPqcjb3k2/9GaTz8u5xEJh7c2oTiFNuWIEYjPQqw74DparUwq
dnVRjKYj8IiyyuXpCtyTgzODA6ycE7sPR+Di1dGHYlulm6VwNDrpH6/byJcCIG9A5671v1Ysl1Hs
oU4hpJ/oxt5aTpuEv4uBJfQknHv35D8Vd7y4TQhglZnPnV93eAnXv+rFPky6e4ooZRkzJPAQmnd7
kDjFT8YOfIn6XjjtOrnxcupoVl4ZEbdrRdeixV7DS9wNZ2wDcBOcbCX5FHigeFcDDRISZgpsF03U
bKZ4RVpOAXkDwfuAQyww2Jog+ghIEYBZKYSfkWRLahjRSyqbafobVbr+7guMMkEmNB0YTF5TtbhB
k7ynY4ABIah80ya8h2lm51n8X0NCAjOQwEX4ab2Z4vzw/KHbDbTKIn6M4tH/Fqtxn5wApg2+Rfiy
orDX9htfzn/zfGv+MKprZjyztTmfY7uAegbTqSXmFlAR5IR4gMpa/g/b68xUPdHgsfBDxM/xuV3M
x0zAzVTmeTHIPslq+5hx4SC3VEFZRVkEL1rN67+P9O57I05EnMj9dnpmdCbN6M7rZaEZvzUiH6Ar
bx+9Jx0o3XLxM36APIuG0r8LC02SXR6dBGC8NfirTnBo1YiWkRViqERnlke9XPdzLs2GYAUMUhgi
D0vnsAQGKczprrvXyodCd0mPKyQ4krxKh7tBAMzI5CgYv5G0+mOPZtAw2bKnCqEDOzonGR6uQgtu
0sUr+CNrvepYls072ex5pzafhbgQsGV7kBZmbhhe2cZCZth+Y4WP0HnTtSFgrwNRVtqqaC4PolBQ
xBhNpoyjqND29Qb0SfhTuEsxxZz5MsuhaWenWMkANeHSaaRX2WDXVhqgxtZUV9aPBzSIJmh2mkAM
1JQ5ZxDffMiduC7hB2//4WAnkG8RSHPaH1eS8AXmfSsL757L8BOyyuYw9aYBGBq5T2ISUEv1Q/u7
SxH43ZRZnFi3f+UhxYKN6wBYcNcFFItAO2xHSYS02R7msKPp8Py+5Ax/PjB5TkY7GqnU7r6TFg7u
Zz7KmrDgKgQfmyizttbeL4rDXzFlz/6R4heDfzjXtlPTr2NrPVamFdK5W+eOuBB31dPZXOK9uL9R
zkw5CutHKOW9owYewbOLJ8f98M5WB9eWHI/KR3pVuTDPfQc594F9Qk7HVu8q+IMKPZakpOv0OlV+
hXknx0SD96qlYcX8jVuLYmX6uYjt8WQMvdiOpcywIeH47LE+dqaGaES1FpV64tCEzmN7Nh25+7QD
74zceK9GJCcKWXqpaXMwmChl2tUe+al8GO0aOyJPIuSsII9NJoa84wjCwoainzBFdnJL1bQ6LZlN
qOvL1K6Q0S1TCurX8KBs4PbA9gPFgSA4PSv3U1EehkL0tJ1QoihaqlTO1TYmuWYY0WU8Iq4QnLgo
JWlkFWhasMgg5qakcThfDCA/nhl71g7S2Bw9zQlsmJBKPs6Q6wiBcRCJJCXHVolk43g4tawJEUn0
39zrxO6sRAuH/H+nsjEGNya3juYfZoR/apVPfHg7ok23pDKSoOgv776bulzXvzcarPVAyPzJMJpl
BjES2WajIwYFSMHdFI4NNVv2CibGkK5H+UzueNOEq5EVnNJkUGOCD4JcT8K2PgxuB1HNIto/0oMg
dJvFhPAosxurh4xdQSuRY4toIKKBEX+76ZfgIXG5UTUoQF33aLj7IrmPrM1yBhpQChWLkUIPdWKs
FmMogOon/zXeHw+IbbN3uNjDQ8x6HW8V/x4wJGxRxJwuFhAjnlbUkCEsnGA4WAoYEZzNfUK3SP6i
YvIdouAdfnA73v2Dix6xXAVSwrCV8dXqgDclsGyjGuw+nbkpvas/C6WIEzqdFHL4+FuWzUIUTbzW
naAtV3p/d9SaET380bheXfNOBp0pbET75d+SEs+6O6OkrPqZFPeavlMA/ciVJA4MdlRTKyQPfr3q
HWhEHbcOHoKRwkIeVsfGkE8Y6CTp1gdbjjmwWMkBGMYVBQAHQAG6mqUkAFWDtQQ8hfOQLz6fvSrs
bicDSn5AvD2D43Zj9hrE+wTZIkJYFGwIGTK8dUdCmLvWF1V9X7hbKRvWAEuO0w069bx1peyWBjdt
8bSOu+aO3uQ0F0KOMuGVo/7bCCERT985l2fL17IjaEc1Wu4nsJCk34Sxw7SxPrT7JABXhA8fwFks
uJDWWAvNTf72tIkqRyv9pnIUXRIlGuVAcAX7QHQ0at/wSUAy/rSUeC3OHXD9LITpd3EX64+f9gMa
Wz4LdaAdfRzEi6K0ObAH3CiKQBBYvmR2Ap63/5NgmRgyjAC3vLK3sY8t3mGAUpcc1fXaR3h1O/vT
2izwl5luUCeih0xpRP2LMkQr4Qy4VzAEDTGHfC9+GzeU4hB3fEOZ4zRRBX7WyIxIifQe+xaGJt6U
MlHK8M51zrnaBnqHsAsCRfJDt3ns0RSiFEsOkF8sR7tcmrLAcqUlhsUJZQwlNHOUt3rG4q2Y0EHI
LG7qmhQsG3T686ZmDfxD3nbLRLdtSIPIEFZCv0/vk2aMwSBFWFRLqcQSh/vdW9F9QCVWU8yxygWt
56cH8y6XmfMTrgoVHnbtk78vbjKnEN1f1EGd7Iouwg5drVJF7aiDDsLBMEXIL2VsO16VMd7FNmQl
zgmFr3yQHrl7S0lIMlQbLE8Ik5W57AbDdrjjf2pwbtlI0ogm7gSvCouXbzrbmNX5F6p95Ha69mQA
mZCXDCAS81Zk6jgrrJGMCAtYacSrp/2xbsxcAsn42CJYpdsq4twXHcZ/T6UeIK8O+mX0qezQEAIo
KZDbaqkCzpYC5XIf0vN2TrMU6koQsma+jPnslAk6XPEfhP9uOXC+eR1Je5nVR9k+f+2esYfyOvFX
Oc1XWehwlH7BiRppqGZ1GKCEeozYANu9yirmVCy7O9E/Lzmjc+x46N78DH4ZwkNp7Qsr2JeDak6F
roIFkcvTkBnlzUKlj/H74pCR0uqmdAJBF3GN89uwcHawPuT3RHH96SFEiuZ5Fhn8fIH2euWo6wd3
jiTvNarnU1BcgMRyUXUx4bW8InJLrJy0xAadPVqJ6k56z8TUhndto3L4zzMPmBt6P/FD+6/Yxf2x
nuF6O2qnn//hffVjrodoz45IKyyYkZw+xCREtKm9Iue2pojvgrL+05v1klurK3NsFGnuUgu8KFFF
55nZ8LnmiwBKMEJhDAEaeBgI8ncbNSX+lOsgBkLxHqbfT7t+qTwsUA2ym1cDxT0shfxPvNmBrwKd
GCMWijGvPkcpD+IwjVMnzDIIdVPWphzkzytlOuFUgLGMCL5G5R9KdkHX83fEucFYqX/0hy3i3mtk
55LbEWch+yKHGGuOvH1HnfAle1U6EnhT7tuEZQawTKbjh1zpUxwmh+rQqGOwnmjIBu984fbZfIqb
+01fpUGFKthRXnN/1pefq2WtzWH2KLAReCJfjVTgRBbaJf89Dnoy0rAqmcpLgLQWuzVXmk9A9p+w
VyCgGZhRxe/05ILtwllAixxHi9BjqBgiX4qc0dRcPo8sYl++cvsyzZtEOvJRsBEKndl0WxqXAqP9
B5tqBcueQnOoJZwr1Ksis3j//ReU3bbmdVl+ICYdj2YDSow/NQOAP31gt42qzNLZNgpEEawPmS+2
3Uz5IX3h4yp98TWUTIEV73MXzEned8Wugo5U8WEk9QzvammNpfOmRfNcEJDcfgl0AsBlwUIV5bvI
nvD3ujmkZ7V+W9rmarlkgwBVm8UqUp+OtJ7WN+cj21QVb14C/K+f82qrvhkWzQlWxx/ASTeQq6TG
raqWFaVc14dahbkD+X0qzQkO42eaFrPb0DeizaBnoMOoiW3fv7VnZTjsIvg6zbR0jZSuR9KfnpNP
ISFNhyawRqct9bMB4SnS2Yc9DASf4E/PME04VQK0Uc5rDBlOvbzhJFgt2/p9w5mawGylHJLzq+lO
ZK4qJmHle6rcZOrH1C1FUEgVGokA4SfqZMB9+f55r4SBQz2AGehwxOYEJqzwKuKNPoytjOegJyFb
l2ub/DoopT9tz5ZHExZXQtzxkvfZX0H2n2lIykdhvh7EQjo0E9vKwb2vLTzpXCoYXTO/pYFuBnyk
oMiXWfgf5OhfCSjMOkI/gYaaurFPX1tP81ulB0D0A0+bLRzFyydKHlvxviawHKNUfFoOIxMsMdYl
eAvMEKbUgg7AL8PIdc4TGPBUXEzIXDwKTzF6IKqS1jcng63G2GkZ+RLoa42v/gF9DIXRAhdqBe0j
1RBPCyqKH9puyQqsHDw4oG5aIVftTshUhBTg0D4o9L+kih8+yMsGywXbHTllyELcLxhNUCf/whP+
Q0PdZ9tSo+vFiApmyJ62Ws9l0w6GdXsOkab/iRE16gE6byli0vll+jtodh0LM4dQxuHf6mx25YEJ
FIwHlA5NQe8ekAWbuwnh+KsVFsYl7t6XIyHq0utKXtv2eV4jKQUzIYBkRL8vwFKL1rptQPXmkazo
jm+9ngDo56XdtiKJywatkrGPoCEz3jlmfETbWjg4plfTB5TGym6vjM1OxeKKP03Lr4H09vWyW1A/
UQgJpgE8oTHZO2SzWmVJDmbQwPQ0bu2o7IbazWwmiZ790J1EwJyQzxxLv2rIb0vTS1PBWOZAB4rM
0LZk2sPv1NKR4Y3i8DMWEG3+X0+t1WRCML0/DaZDJn+D9eFlZVdhe6TxI4iFF8xhzYmRtJdGhcH4
wNXoyEDpbvw+dE3MmPrvK+JhZf1O8JadtHJQWdQ8gUXvvA2PjI1+H6qIP5fixPscCZ0PROtOg70l
q/S8Yo9B/wAw/J/dFnGJjaQ2sPHuebw5C3sfhWlMBNH5cd9dTedZnZRVEGMBo5pnDL6GD6w+rsAz
bbzWwAQNFn/3b3r5/ciVbKLNWSmv+D6MEM+f8Tx1iQpQ8dsxBBTapaxvq39eL68i4uTIAyg87mtr
CVpNmumL/l86xFZuHofxU/n6G20nq53JfN0ZMfHh9bQVn2bO8XkzkOXWpkNMecxyszoSr6m3HjFj
ITkk8i7KdUVLTE7twFpGWOPtZ7m0Z6T7tE4r8990SMLhZB70svcX+fmH9uHKWkfZOh1DZQE6NWkj
Ll8zGOH0zihE44TIoU+LoWULS95yGoPShzVBfkvef47S9nEYtNsbMvZ/J7UL64c5fE2eaXLQOswd
fryncM9HD/Y4iIVL30yTZxEMkeiyobpvBluVnGFF+9GZrizn9rpKN55TVGJemNxbPJOyTGly7Kqf
2X0U/1bstT+Ub++hCyVg7LUvgMkSpEy6ipjAyniq62rZAPksoR1bfsCmTKjXmSLo9Wwk2lAdYVSm
FmKgP2g6wsnrG0eAuq92Rb0EaUiBRIDpLa5kH/qL6p3N5652t4hsUtv6k+mm80GfszCef/rLdGfO
eVfx/IodnoERP/Htp6pXoIcMX3zNY5UTNQ11i0vfhKRmguUlJ31IILPsEaHqa3YgfuJtqOWA164b
VpSvfo5vhCWNQ/ZiXzEIBxGbtxXcmDD2EOMUd0MuoDJtBX/6UWzv0AOtLIchg9nF7btqG7b40YEC
OY7GZCN1bhOHM10QlEEachiuCNgEiNbXgVtPP/GRlJn1+YCyi3uTdhtfAfT2/8eRa/FAHlBT62ZY
x6d6KHFLYZZj8jrKieLmodXLUek+xbgoN8uhDgfKmcBa0YNLMCiaRKGxNmCx1bvkPufwNu/AhOju
4AA/zkQjrWkrF7FvopKOy/+/jmVVvestEUG7rCdcE2rU65Ij/Zt8njA0/fRBew0qcOtAsb5IfDI9
fr+POZO09T5crzYSOELt4NaAKQeRHGT5bpwRWNzVbvdeAXhA0Cp7bgrkKTJdUy68040BW9nQMle3
mHVEZ0K6TTPRMMM/UZKhubo0AX/XYOkl0g5yysFnweZBA0fmveM4XJYV0ym0WbPsvmKQnZMGPliM
TtTA+PnLgpaohNhMN8QPb9L74anbqUW2R4ABL6GZIvVhi/YyJBMIckELqPNnmAhp1X7HxPbIy0Z3
FvOnHuShlHDGqVm93Juf+I0TuAi4V290I22Wi3NwUKMP+P9dRsAISyr5I1RAIZ5+P97fMAG4flgA
RVvTNSBr8FoY7OLbRFhURoOaOmkpRHqbHr4tcZ8NztjEDjM4gKbau5Qlm1nXduT2MjiddVcmgO7s
kClpzFFRvAmhIig+5KYyZEZcZyUwUIAiVz+0dlSGjAUgx57hSQIRpRuZSdGfuh6zjKoyEIZwllSS
j0yWkLtEryW0MzbxNlELyXnEWQKpQOT8PN6zzVTJq8znPQXUf2gKrGJOkxqfsMKukQUmg3Ng8gVw
U1SZahzyLonnwxiXjiMZwNZ/MPMz4937/idm/wnwkvFo12fHf42vNfzc1EVYTy0jUG4yOCnympx/
8Vt59uAV5+RnfU/hMaoVv6XgbNlTsw+/bg86qOiufDhbC2XpfNDMHr6ZWPZnfcBBDlnfXECA2w62
omPKTFneVF1xEqwFZ/kTjSDb0k2yvJ9SWz7qHT1yOBvrFON9JvnVys5adcBl0DZ8wK+vIARaWjfC
ggPPeE40wnOfMV/Fas05aw4L4yVBCGoLEoDFZrr7Em782H9CaBKsd6+QZtaI6SKIyBAJqtjFb07k
zu+1NXT+h+B54Ls95M22U8/kPvJG/TUbHgGwBbl7HtXmoTeHVHT9+UBqxfl4pfRy/cv1q0dlzgof
mphidKvDneY4n4S9tBnut2xkzaPB7Sd6VCKI8Be52MIa/M13y3c80dif3lMCpMru1oTOksXkrnSZ
KItQbFNuqkBibf7CviD5ar/fDk0DRmx4LoOKcQD3w7PssAmgors2/pNFc0gDfPeWAP7OiObSuJ//
w25ZAv+ZyGUPBFrkiSOixfkqhRC3/Iczfq74QRGbuDr7U4//xX0bLQzh9sZa0u5xSgq/DVRtaHpY
ienRB0R5pNlff17yY0ADFsmhGTdzKmQ4oRgpQAMyLGQO2JWQKlOtmxFwW4XWZNlUZ/Hp3O3ipRz+
bRiCurseL4uW1T5M+Btp0ivrdc2qt4r+J4ruuXaCnPI31JfntBO7XZEgbC8a6TEYPdqd+hJf2u2h
cRrQPfl0YFJPW9OiNIEucPs1LedbNSkjCDOApIbwUSXWc0aMXMm99Nn/F2e/5ul/vvVUeK4fJsWh
Gi6AIsR1YLWjmGOx80rcwFsDejL0op5hJwcuk2RlDFDsO8d0e3jYkwsK4/dCUZaqexK5xCuRtBSs
ryXuov+ZSRc8GtuxlOeh/jjE2pois/zeMYBhOf+6aqeLew1olx24VFdGQitr2PNfLkqav7XVqR7s
AWP9eZ2H4auRCAzC5d1g+RlaNbY9IW+cpwk48QROy+9kY4GqLtsJqaqoDeu5wYHanQeXMb8qQ7HG
NEObgnHZPRCIWDcHNt3qO1D5q2gl6TzqsQXVUaeluyaf6tXNzKvUue5DOZc6NfmpwEjqilgS55ry
Z8YQm0uECwaxh5lcc3QwwIdRsKBuUwubdfWmMrV6pmu24blQ0P5wwz1kkuVEaaFCY4Y48AICTF7t
Qt9JqMTnKRVzrQyAc6Vnwh536k9jJZGzWKruZvI3pu8+daG5KUJJ4roCadlWwkavFAtalwOLdZ2B
n5u5OvFw3f5iN2fhR+lYxCJ47vFa2fwY8nyDkXeJ/RcK7zRIhO0muzg935lx0EygAs59WWZ9iV4Y
Ii7njJrZ1HGqYUOpDt6EiWIbwYd81QavFOJso3Fhwuv9+TQhVr2Y1+m9cCz/rFstmgPSMA1gSwhV
fW1a6TEwioSHYSeDsRv59JOpoc+E0dDR0AJ3eOLAgf1E320/ZB17mnqAuz7QVkQp4lBRDtHdbCFF
h2qeG2zICMoY26D6tW0TeXWMAo+zIbSZ5zARLFMpY3rurYaLvTz9kjkxzjOet42RngnegobRrBWP
haxbHRd+cYyQfDvOy2lmwFQFAltRQDjdI5o6/pN1+XXBs6M2rskQChFNbBezCFoGgrQRD9981l9t
21FzKmUrUlfoblAfMOh3DIxOaJIQ5Nt00eyGXriBZTLjcqC0TE7VHhlFrZRKOUl+mEHZhb846nsU
JllwWkROVQa8iSywfcZcPiQG8t+jUjkmAtvbi6wA2tEGo9bnTOc2S/hbHMywc96N5Bt/cvo7+PvU
TPxr5g9pb0AhCWrmceTzDZ09jYGMMVvUmTuLna50saNB/CjQxz0YsbPKoAsoE3mrf9tay9dZ+rBr
pKGHo2ojYgvIRIn7kUreoyBM7sT3ZQA0nXALBCTvLxkeCtrnQwZ3v2+2NBsj12pxD6rBhEY0z5aw
sBoY8WjG5pZiMYMYQPI/Mi5mwkDvIBpE6S4fyGpOIZqypKovl01Vk//BFv8irGiA8URsfz2GVcxJ
QMcUIkRKeLJfiGWEsPlk2Lpfcm1YJ1qWnGlMOjsnOv/eB359+lZuhISI1w/LcF40HFIqagLpfIq0
arBWf2MpypKBADqosYU/kxFvyhPLLcYsoYvA/FHHEQGOB4lKfD5mDy2frj50AMp694fF2VGWPl1L
5AtCIezx2j9+qEQ3QwOsWztdoHblST5Zuld/TXI+dvv1n9wEAmyE6H/vnnDs6ra2Qw80/j0KdsqT
9qQBv59IX3XUyY6q2ky4YecVSM02SdBAUfBjLI+ocnf5Lb+0tmcUhMo/qHz7oGLWDMHq7z4jicOc
9DudIPRLuSxm0qJLATSA0UOC0uJqayxNTNoz5XGD2N4yWD1N6IQC9WrQJdJ5lGAEWtquAPtOUt7V
KkJUJawnR+GjHN+/W1JIi5yb6QSfDKLnWG298ufkTtDefYCIer4Kznf6+mHXQ2WpetWK5NTb56Pc
vPIUBHQ2J8+DZ3AbjbZ/TQzk3/INADk49SXJfhEsxQGGClPy0WwOn4SR+5h0JEbvDf41fPQTcLMB
XH5YQ1woI2G2tboQFkeT+OXJ5qGGYoCrWn9Rlu1mmVJ9eJ5XFROuLu5JwOTiR9y6/3diuy4muPfL
LUVo8R4riYDq3u22kga//CTDvNEtkwd+PoIiDtezxvJjpry9MCx7absLzTF8VR9JvwCuTkH7jQwo
z+M2lS0ODZItMt3wKRVVb2cYhtxvpaLkVwazXDb0a/9BxghQIYxkBoKUOWNszGEpxjyNdZqFOb2A
aFRnJaQmfDxIUmPzZMELWrOLLBGo2iJYwe3w4R4TVZBcy99b/qH1rt4gpNKXpfK7ZrX8F23nG+B6
zj8z4KFU31JdoHRZpnaC5Yko8cbreFhWzyN2xGAyH8aZYO/6pLNLsoTu5P8JhfHOHZaof2XRVrbt
t+oSOqRiWQCa9FLxxxwLUsg4pUdLATmFAxIrr3EDVL/sTpLwzx6HKgH/ijF0TFKWfpgAhEkCaQ45
izeAh34Ueo+es6iwlPobTJ9DWPvK2eDF/sBU5dr6plwB1NRCNpGjeC9hUSdLx4BHDxZGzUhzj+4m
gTxqPDMzv6ymOCdCkHmw7X4y11QYZCDjiJkIaGVaIERq3h75+RGb8E3RBESu0pRO593jIWL9kc2L
GL0NJhVJTPGrcdEXKHgaQ68sz8RDHbLkvW6ApVB7s1X8au3oxe4qIMIl+UJQwWFtNNQhwMSsXFbR
KkcFgyDmXBDxlUpo/maVBE8C35NerPpA3agWIh2N+oY5ERbNURa9sjy15RKqcAK4F8fg2Fonaoan
VSVXm7+Z7p1rC5ldUqetHoVNaSHPgUHsvMw5/Z6ighxXorqCzxmqZ5NaUhA+na3djqvZ8rD5OUrS
9p9gMNrPGHXZ5+gOdgxSZBkmtRbF9L0gcfFV1tne93pfPa/NnacKs8ITpr87zxV9Sa5pGQu/r0h7
WZ4TPbDA2P35Pblm1Q+8IX4pvqqKJoYyScnHWrAHe8sB2XOSp+xUhiKLELKNvxawVmOyhrdRGIkO
JJZrkfXIMiMXFnJRimah8odGRXNK1R/v9zR9YujiTL62lkqJALyFVRLlfcrzGqrl+ZROIcM1gu34
RiYSdLW0LFnWLap3nQ8BTyu4HAfPFMQWyD8970YdLCPj1s4vKyJ1RpBijlxg2mPiA3v/HwBgALnV
Yy+y0KAvm05041j7KXfL2DHdkikADrSS6nUvGUAUUB+Ua3iKuAPvKSxmTsJ22/bUcoF4Jd7Lg94F
md0/3260+QxI+eYQXFrzoRtqiuS9o91IkMgyh5SDQ10sI3u0lvXQVDh7gxzyVz0En6t3s+Rs5c2K
oYDwqOTeGnENDhxTc7anGcyPjT6r8om4jy9esgCta/MYT7ec3xNsnVtLqk3866T84AXS1OvnWDWu
pZ6ZzSzLjviNu0TxhrTIh/SsB/lg91ZH+fuz0O0ylpszX2vdHRsuIet4AKsBbA9j35PuvNZp19fH
x3XhF6W6IlAc2XZym+mGCROSbT2qN/Z9XVt+bcHB/0uTQG8LxPmpq+z1yzT9UEWMRfP68Yh7zOdP
CxYL+Ak3X9CGGRsnXx6JS3Xbnf0JPWuV27PI3gjCOZACyEepEJ9gdCPwNoXt/6b3L3ELS6J4feP8
w5BXCsaup4BB7nQG/UWIQBHN5LFSzSxNLdRsmXpyIUqWYP/cNYwxxZAx6i9D5tE0jomWL7jzWxlY
17h/kGuB/nI/ihw5YkOjqqcSSVvwLJodjO+mLMHR1iSSq/w1UMKaeEFJHhWvMoTu35uvFMECGnUG
IgINVyUeVKppNtXTrS2vrvM5m4Felq3hTiSkbCWjEm/aSNTwlcJclKA4eI0vTnztNZ2DY2H7qIjN
AuI54DaNya9l3oivdZJpDq91RzR3RGQYMx+/1fSz1kpvR3q3BaC7FdIvnYIs5Q/cSf28gMfgi9LZ
Omjl3BRUv+NzD1ARYm8H64/7YaHD7GDhhHBlOWCoLZ7CXk+Rl2nop7MNcCimMmlAGEaTlek4V14h
sSJQKXS/+Q6v9l/e1H1s1t2XZ8DbOD1UilxWAqRH8EJ0EEuq0iVz8z+8ISKmg/KJR4JyD4lxYsFx
0misg8RHs95jURjJPO5Crg4r9dhBQpWI6Lh8ZP2MwRP9VHt3/uEgnpjnmyh7L8aVMTXyBVmE/k5B
epDVVgzAfDivgxisQ8+u5V2ipVrExFNjaVzw5VwNLtNAvkuAtU7fTyfF3LdQBoJUDTZI39KCj53F
zrQNPCCoc+ktxWeLN5sQ/ykJDOOsohPIf/53jJLAQvrC0Vo78cSQ+i7HbqvFvXf/Il9sMl/cXZ69
ctUJfgnemJCg26KRcTCxNzojZZfn1Jtioy2I00LLx52cvZ19P9BQTxqbCrjkD/KHobAoUgVAQkoF
mueDPmO+h2gejp8Hev8OkUSCuLcc35wHoZPIsOK6nymKLfM9lgnUe/9xumzx5MJWGxNcY5r/7VJ+
IHq91ZrIk5mCChOZv+gk0AtPgawzkVpvw4MUHq33tx9cVU3Mi8J6xE69wp7pyIoGB3+MZ9Ii4hcz
Q4JFMNhbzebx/oVxKy59x3pFLmYsH9EGE+w2FYEIsDSV4cEXyindGWcrhvLDhNt0Zy7j5E3oIL6f
trTXuwE8bKMib49aLgzpXWGgYBDK6DBmUTqjQLtNaiVXN4gTgj6A3hiOIQAIshkRwwGrFiVgZwX2
17zyAyEy98DjtkD3u+gafbDs0CpPfLRJaF90CX/TCsypvBVfY7F1p1SNYRUvQMnRP2qnuM4fz6MQ
F5fpJJ65HlluW1un6IcNVavLxNO9/tbxRIjCGPLRsJmKcAJnn6NSQiD+84ximXXPQ8+7a+yV7VVN
PRLt335hkPhZ5p+pbgatZviptsH65HpkBKTdkf4xmnm+1jZs5OeB21BbZyLpNoKdOrNtHl1pdTNN
C/9DwtIgMeR6tkRLl2OE2HJh0WswEb8auPv/TXIBHWEtlw40N7GNp4+8x/27pJSTqahYkwAQjrMT
f04IvccMiIVhxc6ujdsfaLRgi+QHO2nejw4G+QndoiCUBxWY5TKx4inJfAocnEZ0QXCDvubf1Qjd
gHBEudLUlpUJ4az1CYyl8o9+6vYThDMUK+e0V3lyMwzYz2uXxlZKvtI6ow/j4RVUcBLdniE/Nz9I
YPQlKGzvWZAYRwr5qAOMPBvw3WiW3m4QtRRiN+9a3Co1pvWb8y54INgEHNfd+8H9PEGcyX0K2pC1
OzLskVntaklDiFI1DqXVA12PESKpJNa1+11UxJ3vozeUxZPS7fzMrGJ5WifxaG+mIB0M0lnRnXZ6
9ddk9SzFZK7tqJ9ksBUciOZfZGaA1UwiG54xonh+1kH1PV6iXovJ2d6TIch1vXR7YUDug1xbbdGU
tAlZwUL2JWueaFB0KqRV2TWAonXzmywRCE6TTxkVD4V7ovKeaT6GlX8udAtLA5OLBE77lb/LVzTp
ZA6p/3QCw5MDWXiDrYy9kXb/aeSRyWnrawZF26vdXrlqJ99JzSOoV6GuElOsTiDhPCi79mZMqd4N
WVAT0SUl77ClTtGJlgOfO2PQdVpw4dHZMy/nmlcArrwQKY5TJ8M9qA/Mws8wMkv3H7RPbCVQYZ79
V/I4sJ/g7d4O9y1VLailCxJzgXz+b2vWvC2ZSgiK56fJU9uZxuQsrd60PhLDFt518CJUvBf1SiSe
zLNY/FCggwCWA6XZMYcDpAjqyE3i1dGOjfDpkl2kuK4RJZoTNqi5n+06Oalru2/JHYVpgSpU7VIa
F4oMLtOVcURxwNGaAhYCyFrwNDNz8S+35epxYEkE154WvgtcpbBO8oxjMQkFEgNbUWUnlXgCLfDt
e1yrunyq3OJFMrlWlTt9YN3ny8Z+cZAvtrUZQsL/uVS0kIT7gjomsMwR8WjoBrpLIVWm+0u5eFBt
J4jdP8QulL/rS8V4LDjc+6uynQ4BF7olnKFc06WrXLu/nNF1bIQR+qaRFP8+UkENfVE/BqWdyQEB
pWS+EdmATBcO14zwlbMcsitVCIQkAAmBG7NwVLUe+woA0JYNFaiEFtqFV61BFT8q+7impCY8vOTr
hoewENNLcAP0nskMPRkPz/pmRhQsT3Tml3vdFLkYOwvaKJyVLaoL5/H6bl49EuNUqLPIQ5za5nEW
lUCy4CY904q0qvRIyPqgrn5d/8Z5WXS8GVazi83GSwzNuLBri+JAt2lwaJwAQp3XGM/7yV1MWkAy
wXsjk/B+D6gujCIs+z5WDqP7zVaZYKruNG2OllxFptIL3IeeA57p0MRePRoTHxeAuhMiQQ/+YSrY
hNeH+Do1wCrF1KIGU5kdXmWhtNfeKADeR7rWV7g8eO0SrXkAcN9g17VB2knJgE1vIQXAJbEKHv9M
KNDW4KRS0VAHF/dzNwutl70Wy7u8QzZ85m85mpa0Q0DQASmBfIApHIhg+0DbEOaHvBStEoNzU3UH
eTJyXGPpEJdfVrXjft1/Kt6453KpjXfkhLvMixeVr+4VwTNRVcVVCj2YWIrMlRRL5e32P46ASybv
goYV7ubC/fo9mJp8H5O5DAiE3WRwqo3vjqZZIiNvelJDQQeE0HZQaFeZelGLdRU4EZCKmsSEmzhy
Cj69IZhhEGiWqUwaUoMQ66DwpADEF6xOTSzwJnslBViBCg4/+uMt0mq3+MgQY0yqrpTNK3k4x06D
a+tpzk59zHL8DXOiKQUrUkfEkEQ67w96yns8x8UrdUmKg6gqVp+4yTEnOr0GTJU+vb9aJPCxm/Ez
1SMKA2Xk9Sk2KrDkpLJEeXWvCU6Eb5gn9KWB+U8Aay+KbO/MH8MwP0CQcPXpsDn6JIg0f9/L1mKH
kYup76k6293aGhH1PSHOnLbOp+0EYCmFDMB5pWW1NcCqE3KG74fyLdniBxOscOxqeoYM4wUgjBz/
rhGSdK4JkbdrTF0d3to632u5fK0zWpsawT7VaeGvd65jmTSqAqblUfK/MXUFfwMtJ2wapzHKv3z4
T7KW8Bh1QDAebZFE2YlJ1PV0zlWPsGpOf8jRywB/XpJ98U+n41Ti3GGvvuFG7kpQV4+cWHWXoMcQ
8RTENcflrbw4az8YvYjqo5+CNPehhKmdpIs3kHGNTrfEBJzQHXkuNN3Sw25crmF3/rd2p+C/xLab
AZGfnYKOf94QzxVe8fvmoRMSma+aIRsNhG9cnOMuJJ84rAAeFB1uw6oO1w9SRp0KdEG2MrL16qVA
mWjzDGyZhZmsZKxeAx8529R3k0TNavDuubquxGi8uZtQZ+fdlv54uFXXsdSneOtqIJf+DRlONkJw
I3pQech46kLa/HLkVpDL12k8DH3iT/3DLvGJYeQ94+hMOVDIbHPofcWKRwYY2SmChfhCmtZTN9YL
+NaQHRDrHAjZdof2TlPzKfpVGol5Z6q1+DXk9ZgVBxfyocb4zjuHxVBmcH2D5Yjmwwp3Y7rtNxPk
umTp/R45XhGsCKrKFy+UpYRZn8NVdYG81xFbperHksL66jwuC7S3cHhsunYTKAW8sxS+Fpdox4lG
4+rd86SnBLDFjbxkRX1nB4W/Q/3gBTKAdTaFv5/FRFWJUSRvh4Cn+rECPJsVolb7LapafzUWGHSR
4jiFBlSjPWl6yncgg/SJQv10kUo1BfF1t6oW9HcNuAeCrGubMu5mbTMXlHeC9j7PdFZuRUNAfU+E
eqQWX3kJftvlKv+Yh2tj5EIFJLIvp6chkttDhx+cUsk6zh8D/iwT2B1OCDWyn/m3xKcBeESM4715
72e2BpRWBBWItPt4HOo/gem7a4i41Qx3+I7ntxFqH69QFRTwAkBflkWXflmnOHvOKLkR8x5+TZkD
V5Lzn8GBLHzeu5uQ5C4FPH4V94+7mr2K4hnwa3omvioWVtnXD4fU4JnuEzuL/4yx/t4Uhxh19aab
euAjuSyFY1iPh5mWsfP8IYLPUazAXSSE2h37YM0mtJGmJriVC8B6rhin+V8zw0y6h35VbpYqx/Du
l0sDqEiKqWaYIY2uMFJv3gFh/bxnUYA6UWzvRD9AISB4HpR6y6LaDe1jacy7UDjr+oG6vQ1KIvVc
cs2pw1C7b8Fuql4G0quXeuU+EdzQPfX1dhbFEM3G3WcfBGtwyx6qbk4VfXZMxKto7PUAYCoHQTvU
sNLKGU482RlorWoZboubYlumLPkqHa9XxNq3z5WOkZmDP67BLMIwEP9NjAcJU9hbUgNR1JBNBLpl
ofq1aOMPuDqLZIGjLQNZpKHWVaBcY6DA+oDsxOZok+uXtZ5I/wHGSxuchqx4cb1ySwdzxj594R++
9b25eoJHZsI+pCrB3gIgFKpDEiuajvQg+Ewl/A5UHONsVrRrahNMNGs4ejorlH6GmjIwxkdK68Cb
an3/sR82YIk904n2JImypHcMhCFavvn4nPW9kqAvbQqBvtAgu0oIx0EyMeKRf6jzDMECf+YKDhUv
uos+ENWRWWqaW7NboV5dzylm7C+92tpQvSoS0WlNPkKFqneJBX7LAIbjUs3H0YN+rxqaD6p5/DvU
fcHdt0L+E/3nYqxzBeYYbmJh/TPYz9VBw9HUVTd6Rr7qExRHtKikaeqpNqJ63YSdLPuFvmqOLuUg
rs5SqNjtGphwgQZ14bt1PRUca8vFMk0tMaypsKhchqnat/mco2d24RIdqK7+LoIDipJILT7ZZjr1
PQaeQDWvYdN9eVkfWP107M6yGtU1DJQJuz+IXX0slXMZpfHyfFYnmp+ZrPMGwJWIU9BUGG14khbi
51hzt759xLXIqcfhobCFF/RXBiKRXnlzc6b98GW7VVsWgPmICI5SDUFmfjkRNSkYwwZoV8kfbEdc
LB2qEqb0XUFXDNfZ4kAmJWOs6pB4FDawSnRgrflqUgPclZ8yFVj150OAnYQEAK7sK0rIyVoiTuVC
zow3C5Ufo8VFxuLvephmKqcR8U97qJaEixA14ew3yCxG/kM0HZIhPf7i8YTszQupcqfeJoi5I136
Bly9OCLWSUFpTn2lR8BjzGMwhjiEFJccIeyH7DC27BfQlmT5wQ/mG2n6ekHIkVkD8d1LAuLa1Jt1
mfPyUgghUxi0ufnfdU2z2yRUYaI68+uPjSNqNiNJWrKo8BK+GDmKhloJSSQPdZKtgRhgTjjrB0g/
vTii65y2p4/csMlb5l2Jb/SObTv3jRSDuP9/FVbdXmkYiTWFCmMGL26PgbzHF5nRgJPxNib+sFvi
/DXCeoHdvX0Dbe7M2I5tAMV3Fjhq/o86ZUamN/JhqUGqHMliwxmTZsOsNdZMlTsbyAXEZTuF1FJ3
Ri6LoRZgn25Keyz9Cytkyqt62SJT6NzmSCqfvfVcUpdn1dHw4P5n8DPnvhR+OX+yOZGy+TuOTD5x
mDoJcXLTG2ouTtxGEHLQP2v1Haw3ffZVGyJ1i6RmY8uChTOCE+I6/gS2d3QGWeAxtYqn9qaTnWbd
f7ITPJ36jUgYJ9FUwjuWES7iEzTMMzzj9WsR75KgS+5Q5zj17KDexR2QclwE8FhvijQV0KpD8pv/
7UgVLY6fXyH838ijQawkqP7dkePmnNvl3TyPHGuYd9Ahv7iSzRdSvhzOR0J1Pu5g+vX6T77rO0OA
b93rjLO/PvXoMGpV85YZzdRhqCvveoPwp+2x2m2s0+o+1XB9CaGSW7hb+LLT8dnNAMQovCdybfyD
3KOjJifeQTeilhjexODc9oGQ2TSCRc+Ox0u8Wum8RfRKQS2hkt801/+ZVQrXO78FfNb52A8kClJJ
ExYAgS8AC1m4fJ94hnK0ZGIzMOecUzWUxohwxVOqrj7Xx4iNq88zeMR1amWNyaqZvP/KFCes0DnI
CjvIskF+UYXhS3vWGr8AJoEqwhZVR7hozOSEULfau7NQflXQTTIKoJEV2z04lP1ce6Vcf2dMkN0e
kAErI5dA2V6u3b4wbSJFx3fOZ2y3liVanyvfL8Kg+HwcTr7eayPt00z+w6rCw6FsoMNVFRTYhvkf
PW9NmuuwqOLQBhiSLGtaaGun4smcdfcTJxwJEfIysUFQ8W/h0sNjJAkzMk9g2KPvSdjD9a0Bx1AW
lzS5HCEwMTbqi6VplMLYQrdR/Hfs5ca67oAUSLI2IrPcTdEz+7GAIr2EtHGfpPUBraSpoM+4wn2h
iRm2wdebZmtULGQ3+HtTRGUDl5bxrrOK3kgnG9dYliWMoKDW+YCjx2bPArWCLYPGBxiATxUVqOZR
31+Bj1XNwmPx0rMwEoKMxqWU7thQ/9UC+X3r/T+kJxlpp9OlaFFkIvamMRQBAMJOQIfb7It8/hu3
rYheh6nlDgkC1YltH0NVgz0jgai3XjVzFvuq7D2+lECzOMK5oYr+o0azvdzOVZRpQ4fg152x/jq8
ji9jPzpWaNladMnX0OqfaYv2DkM3aNcHp2ibuTm+C8FNn3OELtU2Z3C+8TXADxem009RZMyf1bgy
09Mb1IB4XwLB1/9xLObHc7ID/vb39dksIj09OF+HDxQHH8dfPhrGdmQDGJ+ITHccwl9RdP29G4YY
O4Cwu/E79mGNOV64HnCk5atFENuJuPKn1OzVQkB1XRFg8+hrsEDQrDe/TnmeD7C5zRZADjVFzI2G
NYO3KGF7bDkqG9KaItVzCKN7A+lhxuDSyaouqxgAsN8WUkkW2TECA4LsiOFRmGlVe8ztdt2op3Nx
903GOxwixGwWGSoDwsfHm5ixh5uEm5FYqzz/t4v5zK2bxcYUEfnHEp4Fn1PHhF7MVZVIWhiYbJTh
v1MZsh5xttEZxMupLhXnntvdYqf9O9vCTODA4pGgQqb7RuNWGKDhIPEG46kShsiqXBU3FyET1ze8
bcXf6kx9Lok2fnXXI6Wflm72ji/AYPwMxg4c1TBRvQyB+pHy0WXUv/e1+Bn2qRwyYRSFFy3t/+DJ
82kgh6wFrJbnCmvYFj1q8C4TyTAq4thIqEfXgXV8n5wj83eOz0ka13wQX6GfQGQralsVX488z6jM
s6MM+3srnRVzM9giP0/XT4ZWJIOU4G5in4BZlZ/GiqVWUns5uETW64pRF96zEEX9v6oKME5nw9UJ
tCbwJ1SjiHpFUhaxLB2VyxNtwPFyZ5CeDnZNi2rW1cw2OX8DxRUJEZKWh03PBr4o6MUrCUnXAeG5
EhCP+Cwz/B/0HKNkaucDxGr0HC5P7jwnjD4dbpMEmeWddD752tExw1waVVX5HmJy1gi6mFWIFW+M
Z4zLSE1gcjJ2pUiKcV7s/DzslMQBEIf8m2x5KA2dhRBvR0h/RYAIxuUHqwbJr5v/L0fxBtWYI1WU
RDTRj1x40ZRx99RcgMJ8ZD+eLoEInf2n32l9RCZrLQYnXvvrP50NHvWYCZDYn2bdJ8GjxrAAyfAx
B+fzVtQeDTpSXsnJvEx9AVwDNXE7xwzFe0pEXRKAgnga1n41pnp+bRBwgvsGbstMtI8e9aw7Z+T2
1pnAuhtZEGVv+TkSxcAIQ3SSKF4PxGU5Cype+uCk0n+b4xdHECvVIiSyPoZ1ZepnurZM1gRfh7/Q
wpMxmgt6zwUOn+dZ2TIyfRfbmGDgdLXnR69YAPoGxzpRlD0WOWvqwyLs74vs4McDS5u6kNPxKJRE
SG7Z9k2Q6UaY0quNf5yC2NVx0KfGSLpqSsJE0TaQRq7hO6w6VZwPCcnXH/yv6IZCuOziyiQ/8rfD
LbAl8eBYmt77DmYe1uqMDN0KuotCJkPFs+jYPO0F6FW3EtAlBOAGYa/lbRIUwiEj2AfpXPFHLCz2
cOlUiu7fxcDiYKA0pDh7PW7UXBrVY9x3bBGM1MAUMVLkWXf9CbiWN0+ZyXztOLqbULuM5qytBp+L
QKFHfdoFpXXnTR2pPUf9wv9l98urUA7CqKxttZLXklap0h1vVgGtF+Jo72Kgx6Vw70Emi8bT22bL
FJVRfKPUO81gXa4BQ/Y/noC/l93Q3K5dymtUOpcTQ5F6pnvB1vIOyNwXWYlhZvHeJsHO47LXmQTQ
trZF3PzT8j20zqCWAPgfyRJ9EWABtVYG5x9xy6Vpg2jj8rmcdHmx0iwwx3abmTz3cuLVaQ2G8a3B
mmFLiy4K8RmSthtqAuH39XMEgD5LADwfT/xfoFKbe3HBcDcq+PEGzOODTrwZGfhKI/2B5Jhfm+rN
w2YybMOjj/Brrim9WkXd7CZSlIkbc8qMlA7r+Mx+psgZxFyLnV7sA5U09SmqiWXTPjt+0hfW9Wcn
tFEwugqjFeVXgululZsn9obFNlMImnmh7lmngBInsb6ewwHnk1jmQsapueC/R8Hh7uwnmoHyIYcI
31ahiGIfJZmFEuBhILRT8PAzxP4nAheNEWtR9uC+k0k1W04/JfW7D8TA35p1l5Epdy0PO4SR8SSy
w5nl0ro2wVIhriTkQXZjAt/ewn1adwZrZeVIt4zaKmOyKZqo+QnO0jiEixL4bivpTbyz1hy7OuCW
IqFc7Lk7A9fKoE5VjEcBfk6b2z1Yf/TODgaloBlf34A0yxkTI1W6Qp9gMZGYpO0SSjsFCR1R5t7i
lB+12wRI6FkB9dkHA7LRn6J4uBmUMm/90aZYFGPE5AL380PdzTSrMA5fHgM0nIkKidNRZBuYlkC+
2di6t5sUib5xAQ2ecmJ9sEKEUF905qZPSzPX1VugJzQsOA68qXCfwqsXdViicfkGImYjbb8N/i9Q
yOnTWxy6hlflZaWSZFbHhmuwWzcOuP7cp6dpzPy18KhTH4WlAdYuFicILPe4jSSLxrzpy6NZAA90
t8xtuhRhxUpiwL0U0pZzAVdYltOS3gl8BnzBeadVnFLBq6s0MpHdPTr2pdYlEXvDXTnTzolJl58o
lzliRubPyLTUt2luPnLFRTluAVLQNmrIObo/iRdEU3ibmIY4DL1QJBvuigW8IwBXxo+QpC5jk4R5
5bQFrPfxff8Lbmj25ZNy35s1jtppkf95is0vSjIJhR75Z0soOp2b62NG12EI/tKAcEu5YcUhMAiy
+9H+XEiRgfNLiN8pPEeWN4M5TsP4HLUlNtLycOR77i1WgY7bLpq3oHBFOGw/Th1DSnwMx+Qdu3TX
4kk+uhQNh+T/0277hAa/b7RYLTbT2gdLuzIGI4207vnK0fZjAiQnaOmBAG0EWPqz2STWVGOw3T2W
EFtrdxUHsODnYXrgK9N6bQdT13p7RjXbpujG2PJXGiJGhtuhxllqN/Ml2S3BUKI10dNM7R3nxRyR
C66zmEoYM8KEG+gna/212jq5W1WEIni7X7fEPJzlmKX0WLoQ9WAUmHv6fagP7VRGuPnsdvHgEhG8
d4OTvV8kWx0A7e6ku/+95FD3kURwzLp1NtXpsc0wE37RIMsdVGIk6aN9l3iWlXhgNZhBiOdNiyPk
0C72E44eeYI/UjrncCTSIViUhv6Lluy7U47CMVI/6X/4IGLQ0y09u0mAB9IzaLgxxZWY5LzaZjFe
glASv5ZA4475PHGtL8Pq9oVD1N5AGH27QWo0AFkbD4ifUB5ThDYvB4Hwxru3SS3+t2/2Ywhhi2k5
KmX6hBGkgu9IO3ByvyGC68C2+ItBj27L6Hqx1bQnLYgXDby5N4MJqda5LeVAjhGW+N4jYDalrcU5
on0ankdNLuIsQwKi+zJd1aDzCq3fQF2Mf5BRI9xGQDXcd2tGLvF5J/I9gbrRruSiEp6660arJ4Qp
KrJBYzF0sM6aJ2vrk4Um5RaMOcyyVFznwLABUK9jJ5AeHtkp8YqAuvHEJ1mpLbmOzeE0y1tnf9Zi
w2I5RHa+Zjrvkh3cy9Au8qez7FjmzqvoUlwnU9H92HNHVIhGS/a4DEddaENdJK9/gXqRjQ44abxP
57dv+DftaD1MYz8Nr6hEyHwRLoBp9bEHq6AKoJiGw/EGg3Heh/UwbE0vGMULZT7D71P1zs7G2u1Y
PvQraWWuG/oURK4mLm4l92wH0AKR7dr0l1c6OoXaTaunFPtErTwIBqYHLl26G5CCuAzprsbCgfzA
cgFH9av5sliAAk2is3yLR2oocESZ+c6aU6qPKTSs6ZPqOojyZMX2bLKXpeVhZkSTV0tCzM9UmtpA
G8PrTdDAcukiwpvajBv3hCpyfnKOGxxMlechlfbN0dMlUFUZWMVy6EC9xqObIXFmyZyeVYCGl/LD
caq3PFbzboJ5wLHXOJO2BCFDucMhP8R1IXuZEyupeO1l46qKIoPrhwA8LeNtd+7kwcKQNeXEgWjE
lh6kLjUMtINaWD4riklqxC5yo7RhxQJLKBLqS/ClSg4S65tv/znY8rP/w7mFALKboQkSx5ZmNFss
0yP7aJID4XHPKWCWF9vhg/YiZa+LFrAfj9TpelQfYzkcwTq+9Qaulwp15eKojnDBR4yzZDg5Ar2G
sGNUSquh6sldpTDNGGxsDCLasFYxiPXe6zZFR2m5la4CUaPUo1lpFc6PHo7w8HXhayM3wES3vmXp
jC9e1uYF70Sok8gMVyGrCfwztiJzVgRI9EMRbXL8lA8s9ZHJay40q7k7ynGYpNn85MrJGEtYJEDf
g0IU9ol3bdOpd34cjfdpMJj7uONFyhTPgvJ+qK97ozH/X7Xxgdtw4SDpfye82TgZpy+DfUScS/9r
yWcJjfjWuGDZ97vMWfcqGO8m9jfpToAzcAC8gumds9BkoBy97+Mxn4Xt0prY1S0smVkLtq/mpH3y
iVSxa3HGcmR7nHoDVX4prtxL1z2V2Je3+P+GZ2mbW/TKfT5sYzT4Hy0ZEvC/vBhtOyle3Jzx7WXN
OFt9et5dRYKI7VwBABLqYXCteUanJ6+Rxs+zfVu47NXRz7EYZDdND6q3hzh8aXBmYdGusw56hqBo
LpUtOq6QMuWmaPQQksjcNUBnYjIYmJltPq+4utFSvw7n4fu6fWntgDzNRxixORb/e2hgyl0sZWTL
o2obsC5Nut4Nz0iG9wKqqAOluR4p8E0bDMJxnJXhWZi9RtUQUQGgSBmJX4A1HIeY/wHrO/ZWKBg1
11mxUJUtRbS9HpGVJOkba6ZFf6flS53ytecIBLF1hqVjwXRcU5qxpui9mqaWsgk/w9rs+WRnDIbi
v4e1Y1jj19AzoNARI+sAHYbR/dw/IStl4sTuUguZoMmV53KtmgXZlK0c8LoyC9T9nOMQ3uHRv6yh
5lrKiza7IGD+rCJWRkf/K1O6mrYqCLJjZL0OQcVT5RNYK8I8T5NoL4rGEUfPoGWbV9Cw4NigDDqY
zi0dTTSnAq2eZBGHeR9I+O07g3d46hRkpAwmu1u+n9lNX7WJdgT7ZNubxFUdB5vqXwq2D6Crakj1
zwczLQUJ0zvZsvMrc3b30rTWrEDrlhAVORiB0OioCVio2LbUirnsjdwMdB+tnNr1DSsnu9zGoK7s
Ooa43wDX4f6uBNRsbhNRnQ5zyr0zpO6SHyY99wDeEZoSHcwtIb2k34x9pc0Q3nUQ1sySuHGLds8j
7qbxwXk4bfFPj/rumR5BWFd68h/xb1J6nNDsMgwlwZHkcLhgqCG3P1EFyxp9pdqnAR59L56a/fzP
1zb24gw5kH9wGLo3wPQIZ/OQI9a/QtCVBRIls6jOM+OTchao+llSm1vhhhGQ2yAw/Gqx4t1geijp
xvcGdqw4PkqqPjEvI6QbJtrmz+khlKa3A/ahNGVY6/si7ByZ3g6KIE15VgruS8y7pX5ClYkKXvBE
IUaEFEmpx0WEHfu4nbp2FOgmw49BK/kvP2ff1yOP2RJTuqz0047NJuEFxPsZdxnP45//ezQ8Wopg
oJhlg9JplpbNF28uaPiqZWMJZxJ35u3xkBTPWY+bpB6PCfvdKw5+PhpzLa2W9ocb8Ky7a2ID+Cgj
eERwI9JwIbznl/SRc4rOzH4HV04QQ5hbw+h5H9vgvIQ7Csh1ty8sir4FnYIxSsJAYNZarS3Wo4Ww
MAJwOZ4tSirjyn2TMaSWOz8GaxhfL8m7S7GcUcEzbbyckwJ6hNIZPifwscTAPKtSzx9kmcqCxrUe
idT6FXbVFaD8uciQoguTBuuPrWMFNINnIcq3pcyYWpg7bt4ZhEXlZS6NPNjJ+mYCi2mQTCL85mSt
0bgyiNYXoOc/mXGcnIJcZTo7epZuunBa0ezsNGQcS4wVVVZ+hvSCYSww+pWiXw4vQTEnAttD3Mcd
gZUiqCOznMb9zbHxx+Xi6LfWRCOCoGkBgDaXpMtbQMasol+ltIlZzrh//jIS+b+03gyhvMDdxp/n
Tu/1ztwSn1/bIk1OXGehFFJ+dr0fHqyuXbxOKfcYxi3ok6nBZk2Fb6ahMR5RiW4SzL5CEckoYgUy
+VpZVPKoO4O6WPs0+ky8UY3HUggiEep7npQm/G/aYUcc17bblNwX0GC7YDn9shHugMFQ1tHkg924
8zl4fQzk56RFgSPyLsf/sJZEb5Jl5OS4SGjqqFUEiXdtDaXO/PJGxb/JtF83Xek7PBrJU31Zfr7N
Yw/THJDrZ6RQOzIJ+Z3RnYaA8FQGndSUGlBcASIetg3KsLcpMKpgN7Sje9N0yZ2EtNAORncq2/qH
Z5dd1EyjP0JbEbxDYHmtbleae81v6CYprj9snUDE7HiMcIQ6juhusMbb6vwrUPx6up7pZMvkZNTB
wEHKqXwwveSBjavBZxYqOcsg6RG379XxD44gQWeS9UqydyDGgyRMmwjfv27aagpY2KC8TQhZgpM7
esmbPUyhZMHzBWgijIaNkqhWBMUhi0U2pNdF54FbVbKly/VDQDZs+7qhrPRippOML9CRXBKYGGaI
uD7nxYcSbtWwCJqFPUJRj9r9sXGjvX7A2vb6nI0UX0NeI2zB41eZkIDOC5AQF/9t1iWJBwAV9g9B
gOQWUt7ORlk0TeiFnUA8MKHvzwO21SazVfJm05lMZeWOd4DFjRUDDEFN7NlosR0/Ni2naFXity6P
Iu97X43+dE5qnEfDq1jQnISdnPAzEt7MwzGTPhlxJAyRO//vV1mHgai9Ft0kt/vbUnWfTFGtWGr8
VAW+8IlIF6bawDZ9jTH5uG13pxROpxZSrjgwRApHeWhK4rO2RPsmDjj3LmwVpCD+O9SxXJGvEbxE
87A6YOl7z329a4b3MuwsEc7E+w6r68325YJ4rFhSaDSqdEJiI/Tsepj8yBEUDQRmSpHmVJ6N78jk
MNRF7M/gSgz2r0plWXQL0DDO9NicbtRGlsFo+eXnLFvPU6tRr+PDszwXQTs2D6Ideas7InZk+NXJ
1EG+cvWPUu1gMYO1mTQSIQcHc9LkxjVOKDGWb9s+nWE1CkMNMeysko+OW2RfcUVzCCDf5FFK9UbI
R4Lv3h84cwXw0SrWpzlT4ctAgmkq0FT4nVvKbQckQBBdBoUu1+rGAJbcmonwWwR1S8u8HChhk/S7
g5cDhUbodp8ZMsDo/S+ldd0T2flNgN87YIOJxhfmGoUWT+J2WYEHyu8H/DWjnb5v/bLc/qCvsK3p
5IAoR4xy+wMpErevqXpfMgPAm3M73XDgUdLtrmhQXCua2B7fHrAc67q9qBHlT4lWmHxO015V8auE
FTLqzV0B+tVYqSQvKpmmKhh1sXF9nLkWg3gs0ryik5B0bRn3h9lF/tqlmU9PPhvkNQ9GaCWsBiFi
fLUP9G8wn94L/OSp+od1D3hwIwAEgu/izpx4g6189+bjGPhq6T3BSukJd0SjHdy5DZSaStyox+/b
Jd3eJjHM/+HA2TSSb3zTyShnjtwhazRiifeTVAQmjg9YEdzg3Xo6AGeBgPH0A6dp6G/+dgOAonuj
cpt5Kv0/1rUL1LcosTnjqUqR4dKBl0DB+/b5RQeZi1tRPtjQZBC2FbNly3I7SzKyGopmB9rreIhy
l5JsOpIjlJbaQNPNQbPSKOysarNBCbTK7KYnybaQUN9aPgURx4wPvP4Jx/YBIeEkFfVObEvw6Kme
WTIDwN1Zku7ukGmWzJaW1YsTmc6kGZzV7sjBMPt536TtFO0zxPSiza7R9vPO+BnGPbYam8nbohGh
h+W4AXeDmqXw7/4tWDctg9t6R4O+hwMOaXx7mS3UkMZYdnFNy+1oRHMOqK3yEDiLHLgZJkArQ+96
WtL7BxZ9pccaeoDmIUEX8awnwRmKg+MsKeE9PH8z2QDY/F7U7UvyZR+Yqy7iAbDKs1w2iPuQHfkQ
N1j+mcU+lK8zU3l62BbYtWSzKYcxJq9we3CAmdNWIOtFSdJzMAIYRpCJ/S7POicKZCJsCjh6m4qk
ORCFBqKnfEs2Fsk22M5bqHrv52rcNWquAaZxkng4cxCzjHpM2+Vx3LY99XlEXXsT2aUIGpHjtsLW
y/1mfBbyKRXtHuqE1nPWyOp6SWnpEH6bWOt9X+ix8oPz6phEWqKfuE9lzQHtCmK+C8I5tIMoZQLj
XGzxLCNtm2edX3IhrWC5rvCohY1pzP7EiMv3ZrpTUybx0Z9i3H9Ki/CqXHe6CjPB1dpkf6xOEY9e
1BC00JMn36eikfHAsBQvO1vhCFDqOOOvQHm2R3MeGU5DiIe2d/anduXwo/XvncwQhsRYbYQ/MwD3
poQFNRqmUGOd93SHAzLQeLZbjltSdj1/07GZQKpl3uIDUWqZ4EmmnpooA2NIkxo4HrWCOT6HUuPf
va8+N3xXqmtQ8HzyUG9IQb9d2ToqK5tDj/FjW1xEGGX6fAMCGBZrXu80g7Y0Ya2yo7+vyBstVv4k
hkhCf+pamLEhCbvvktbCz0yDZ48TxlknpCif/0KQtAGZc9qMKCMrJL9VErAo3g2E2PrgLB9XuESU
1oRBTmkT6offGeUoldVlXwIycuMFPrNaj2IPMTgR72qd+Gy7RX5bPCUXwmF44TXXE3NLil/85zRH
nAZaUY4r7v0HYxI3TK5RHZrvYxJE3+r5nUepHqD167gvdiDnGBRfuATCFepyoAdedBa8ca5C4SVC
bbvQP+fSezX67NiuzEcuF3bGgq9ePdWoAk3ixqJQXsNjDMBlfpMqXq7DDiD8ouRYBYVhdWPNS0Lj
XxmIxoJYs5VQJGlDyatUCg0HORKdlTHvLzmCeO1RrcHg+yAw5LomjIIqhs65yUqVOfklRmQ7Z0vf
my/zb7M0mPd447PtfEYmPc93evztLJ+pS61eYH3+7ayqf/7mJixOQ/Mnf8XaJ8d1YSZMYgMWK5e9
zIkbmXd+OC2q4mtLtFQ/byGHBkNQHa+7UMuy9rDNSMCRFemurrjjQYlp/dXLZEqM30p5JIXijnCH
5ZbazFBRggwR6QVx4eZtvRGQL3KC2WTJ7eBPYIQaw3ZuC9dO+Zzygl/Q7Yn71Fv7WPF4Z/AA5v1R
OuoKwpkqgZnBiXk76jdwb50k4KwLQ1wPOOwLPKNuRFMSs6RlcopFYLKScPFd3KejuZNRMRg/PUvI
1Zz0eNl8z3mQN1sNwj0YTINC7ERIXucCRKLAXJKHHYbmIkjvutsWUOn2Fnc9eS323nFiL+9m6+Tr
9MUdkRa83LUHxvaQjAqOZOvoz0EAGD9E9ADTkNpjmja0hHWeRC0OsTHeGNmJ9noQIKUapD3RxrUJ
3hvsGOgHKyIrU6yxbUOTxSd6j2bJSd66REQRVxfVJVArycp8nUwatY4WvkGeVqe/Zo4ndVTeD6gR
DLPxYaKvRBeaB4PnacGdtfT3adAFPIigTVHiFezE8zew30QW6qy7b4HrHIbT2Ldshe/c77L7TRd0
h5ps3+su8lJCFWR3Mi1xCyMIrXXgbcIzXTNEHltgcIfoXgKSkNCDVpd/JAZpqHkvH4CVIo6QcPmK
h7bSIrF3SrTYFnQSQNxwCucBj3HCk/wWjn+61v2d9uNWGll89nseK7PDGLjQISHltnKEYC7WpJ2P
avmC45Oh5ems02IFHR4ef3Slhb2qG3EQ5wRtAmKEGja8KYQKjloEZOI6xYD9ti01Df+RcdKePA90
e6eQkdsRpqA+Gfx5YNi6OttitnlGqkX8VnEGpaN4NqbeWJTrh4cnzJpau3nVtheSPJTS3qPRFKyw
t0YwxJrTrpmOxxdCJR5snecYZ75u7GZRVhUKBRt6Ku3kpoVdIFnIueqMVI44yyW9YKEjBQVC9fLU
JTPj49X2ZPFpKdGDsUU8W5AG3gRhR+JV0/tJEbWz3S1M9j7q1Ud7k/SIw4mBjYfuMe4Bkk9WvmJi
d9c7EG6hLJ41vmuG/9H2JS6AkJ8U0XG05Hn7+4WXJ4QONoWdds7kjhV7llac5l8W5i0RguC/ZhVl
i7Foou5KUprmFHN09RBazP3A+BSCgB4fhPzwF3H+9K/mUN+c7woVAH4E2zAS/8aJnO3pT7fq9qLd
NpsiSOBEuC0FntH53YzpTTXS+c339qJ4ZLVVGuaLDa2CVj8XmmDPCMrzxmwaBtG3ANaLHQM9sYuf
Myeugezv1iMhQlgrRzru+1YRGCsDRNGk230ZpPcBj+4vv2Wa0U4JnKQYppmEWUbREKm5Pppf5ZA8
M37REhE5tIE17xh0w8AOI47hDro2Rcb549q9gxoomC3FpiLFLkaAVMwOb3HeKcBXIZdw5Y49U8VT
3J9PS3w+l2RXi/zZIewicDWKiPCTSjdogGbbkpgEer/G3tOA7VvfpOQ+z8h2H6oPB4yYuXSlezKU
HhmeKW28E9js0VOfh0IKp64yKJG7Ak1y3c9a4LT2at44We7nidbUyAOtSJQssJxGkdwPiVTvpRfA
joDzr+Yjwsp8wRGizGP0o9dTlieRQ2Y6LObIix+ZMtv0y5CmBo5cdhy9QuYgsk7TQynD1prqWLs2
/O7CUWjuEGOgxi19CUEOoiII8+D/yks5ju2W9ZALnonEu506C9ZOqCiSL0v6SJv6ouKiPAVp8w1l
A3JxTn5SDKVMShHFQncsvCE7hqwZYZNStSbo/n4Wl+RQpzv6FSCW/BFAH1AboM4MEXYBkPYi30/I
jXS2mwPmSU0eFR7UaxD1DS40334s3lx6WemVJvQMjosmSgxFoIb9x5bqoNWU4uZS/FDaZL8oBTFb
CcWbkqtRYvuPLVzMGs0aoLjY5Gum6dTJzMIZCO7VAtP2X0s2MzWiPwMRWtrDWo4d02KnBm9jBeHJ
OaTQaPPcuUpZi9V+5NxvHZAB2iGuY5G5jzdYIo9cwvC2+X3jUU8/v5GC8BeaaZVWP6Z42qyrAqPN
pSzHaJ7EqtfLXqg+AvrCYBTcRfQgyrCDpqlF/L7wMCJHqiVT7vH0ns2asVWsKv+ijQR0LT8jvXAc
odfXZeie4FlBNPfyGZEn48XneD/oIEi7oLWVLFFzbcEJc79cWufhUZL4C8Ng/ZzDd+zN1+xup3de
/MJkuTr/J9Rr4/y259zTFVkS+3c4rz0KbzR3UMnU9whc2KfkanmZVweQABWwXJ8HH6/Wa7UUVLJZ
NslpACbCOYnN27cHInzcQgO34SzQPJtKmtG4Gr0HyjSBaQ/XxF3riV00AszNui3X6pgxXqXm57jF
3kykB9ynrzbKPvwbwSV/TD+h7YtOJZv+ZeXv9zwMTRPKZFoRqNTFnTbKT9Mvrh1H8HUgREwD3mRf
rB+B1+fXklbkaCidWgpArbQiTUfDAUTIJiX1wUsIMQfsyRn5LJlThcOeei15A+mrDZLl/StlJycg
tKZrva9YvMMncu/yk8S5CzVTItxbQlWztH8mO+ySn3g9KX186ikCA+fsJLWmIfImI5+Bw4LjEEnr
nsmvvrCZvhc3rI7Uh9PY4Rqkj9I8D7v3FDcpaIxBK4mudIyGSCEIJvxk+g3ezqvb5SOYuJqfm4D9
MVQFBH7Uqa57retApRun4NPxXGyJkMo2gzOtQG4IG6I5Qhja9SrGU0yaLzSTIwmeqvEuIa/Q6O5/
ogr6M+r840vNumR0NOJK3F+G61Oxp/yMhoLJc3NCICcb9rgAcSJHjc23dat/pXxCDKk7aR/mcBWM
XDRZ9wDlvXY/B6h2p6VAAb33fuaOOi3JWI4HqZPHtHvsZW/2uGludj8Ynufas/BKevwMY9ld4MWV
fDSswL+SU38J6fsbAq2/90z4UrVJVpmLUCFpy4GwgccsmZOwGVP+TGDdMQDYTrWtBmiXb2mvb6D/
vqBK1KJSVGZSO57LItiPJbfsOdz1XjiihkY3F/tapXC5i/bbrON5cgfmVEQoTI/SeE/2RE+iJ3Uz
srL9dOYwAbjjR5sx66WtW29wAzuLOq4DLkNl4rkQSDluAJsMjTmMCLtRikqStI3pwDuKVmgixqGD
NyDxJ5VhfE2uNlvagdhJPkVTeGtqhE/4mJ8QGlW+MK9GCcymtJOjvjdcSBl7QnRMiQ5j1qQoP2Ms
ZBxY+ACxyAl96Pi1RuO/fDMXupk0HBgPDFgxj0KbfMikzc4TME9xYf20LlRA0qcfWqvMsohkmKxZ
+cMQISU2+eTz21K6FjdBw9hIBCstw6ucJkGTX0epNRzjvswBqEWwnqXFLrgdjOi9rO1qjTCLMvls
qUfJgf5XjGivx7jvcfBy1Vf3J+qhuFZqhcKGNuqHbnxrAA1OynvNs+/PcMnfGTmg5734AkbQcVzc
sO8h2iueHsjroiyNvxeytXQk0gzSczDdxMuV6YHmJ42ndcQNUN5RrPTEA2lCNYaor4Z0RltbnuMM
WNG7VaER+fpJSYbkC3DAIAWw/NZL4LfVoWAZO8WfW5/HhuU8Mp4Fu4Zc0O1fym5APj43c5exaRLZ
gY6goz0x8M6Rp85xqZFEPX+qOrls3qqHXWuj4iULrDPOIQjfDher3nxveEZDMgooRClKbAZdy84e
E/7fmFaCJAdXyCx1mX8ZjU/gIlMxqobAKYSiP4P9PAlHOyYuOQk11jMOEERB4ta7ECHuPCJfDDNg
IL+hUZttPuRrKgCC4oC2DcSi86HJLlillu6dgOzcIlNq9BlPa/YIxTKA9ZkvN5o8hp93cJBD6Lw7
5R2FsOuCU6TWy1FBmauJalftS1fLBj1H510/ojt15kIGUMHSC0QIZW9/8bpULjggJsvxbG8Ik/1X
70ICwf2On3C6brXNOzIxqQf65LKiIlbluB6sqeni572oLfYFViuX2VkDrBcdkJPdaVwwgo83xNK/
2kFmXC5+wOqnvZpH3ZWxukWAvxAkSZHDsf3UbiXfTaU6QF1oAhH/BEJUG2bcIHHjydIPj2r1Tvwm
5kWDv2DzzGTF22wMFQe3e1u7zRyXyaTQSSHZa2lCGcAVwZ5k9jGhtRlMXTiihjDXyxxYgfwhOkmE
ro/Y2V1+UdNESIT7gmFtMxfdOOaTEiudp95jwjPcqITrPTPR62sRAwm0+zC9A2T6H4IR0nSGg99d
LsYJzbesEBUeV7hT6OJTe1hlczRuPb4IJtH/3NqyOZQm4DR2UlKCfgonj8kc2ctgsh2/XJQRgXLb
CwKydNi9wqfe5gcmcnaH7tJXx0Wh3RV9SYiL7j8M6Nvh+jEVdZ2sCop0i7wS76gu8jcIrhAmsTT2
v984ozCOJ9joeuhh5m9Wsa1JW3U7VIIo5INUm2dR97uygOyVug/CCJ+HU25f+kLbHwyGq8BsMLQi
BHtfsilyfNhalW+AsvaHHRu57dHwC+FI7jNvCGEM0qTu3tM2RdqQRuHpLcEeqxxyDPn9H4f1iZp9
EMyTZkASXZygdxmHgPxxRT1vAtKuWqHmqMr5+0SEfoOP9d4Pfg1M/9lrMhTGZhgkLQWPfWNRgMEi
zTXlBISyNbIVS4QPsVWm0TFV/H1KKdy154qgiNrNXjFXH/G53mYyHDXNyQEf3hzhrJYy/NLB2k3c
GVArKbm3yu86gQnpC1PZj+qoS/Qocg6f0WfFR+IcS6RIRTEoMwYH6/cPE5mbrLZNjR/+fs5elQ9T
x5yB0Y72PA5k6nKbEjYWHO0fGpqlze2a+pMt8NgwZsF/4PczUJY9mVK4x3n3kr8MJW4XQQLtTydU
hz3BEmH5K6Cokrd1McyxmjL3bWKO5J67VWFoG/V+qAp+DVPCFxwRR1d12B7ob1v5RsTW0t15fYMG
SwrI7r0fNwrWXV/MRbSAFtXKr80K1xgORWEM1DpFo+D2yvZW3CH8J/aLA56rylyAUtZCWoBg6rHV
XooOrAl8mzP9FUuyspeWNrCyL9sqwv7IWLi+zVpDXdozXSlteLZYRwhf106Nv0PgqWrceBBz/K6L
kL38ywizeHUvZYTj+s5D3DC6m416jvlXnIVUrMTEzrFXPywMz7LCy4nEpryP2KIK1hyC6uK/mjXC
klAkCZCvXi9ZyUmSoEkMGwO8kxzLB8D9wCdtzycnCu51Yl0dRhJXMmSbjy91T+31FVibez37PYiT
mFL+q061ilr1bvvZHBebdBc8xuFPbLuesYbnH9orqFLKA7cQYnNZri4O8mghThAdOMUan5oSD2/8
r0jntu+0r8Nru7YEmhgU6fHtnkQ99XJJZQfApXtwA2clmAh4tzYHFgZ0BQg78jF4WfDS22PAFaG9
HKvqrPbm1LCiFjli/PZeoiAhAX4rrfwV2hGfjsFDhCwgW+58iAEvq1QrQsr0Awkj3JnlyPZEEbK7
XjHS4jM4TjSMOTHby7wB7+r88juhbwc+bbkMT6STtaQbDCt9UKBbYxSjM8Y6gpbaBT39v4TjHYN2
clyOL4vn27Sp3IFr8vLHalrIDm7f6dU6AUFT4gh2YCzCSsT+8CEUpH8aHoSVGOgvcjZAK7SQJ8Go
/SdfwtPoKskbHhHOGhSmkVXh/XI/74/s1WZ3HujvO+0QXwqacRTfyVXBhYiya6kqeDlUqNKbElGa
nhiKLdhduGZcjo8Jx8vCGXg9mcxbLF/rZQyupwBgr1g30WWUQBoDRjOHpq9UXoGaspjMAUj6ew+b
OpCeOfEblcqtaqMzZnB6kTmTtyDmLI/jmaG24Hnx62gw9+wsnO3PTCnrnzXNpIS2/JUd4s6Lv5Zi
iKwrjebXCwGu0Vwabz8gHAodprO0Z8eCf3UPyMJV/9qC227ytn3HQze8U0tVy3pxoUWMmJcnEIb5
6xm2rimRy/58fR7beOeVftONc6ajv1aKiQeS6EGGqcE43xAtEM9DP8AiKhO0Q2pJcr7zj0RVL77S
H2GJ/C5SkMLK1bPW/RvV7QguZDweRNF3+bjl38dY0s7+2wapZoE7AIrP0+bxCu21V7XgBT7Jj7FZ
LS2Iooc2rQiiDQuQFmKfH0/2k1b7t7QoDfofC6jyfc8HZZSkN3DqMCfVj32q/5IY6U6E1EL3Ocgk
HSx/Buig5b2YXwRjSEMGz73kkLHKsbnBWqjUjIP0c6csZmjv6/281v2+JFdtcX07PVx/yQf3czay
aNSSjDuja0Zb8D5Kpq1lTEqqNqkuTK0OjIgsjlH2iJTjgweSFh8a/0A7hffO57mTLB0Jm9zAhkrR
KrvRF/qtg04LrAwIEc3+/C7tbvufj+KCdx9WFe9sFYbqHoM4ULxQgZWI9ePi2qeu6sFxIWQ3d2uL
ZQGjcfWQReBGotsLhxpVgvy1QJEiso0VAWYLPvTiY6PpX0GjZnO2ii35UHaS3oTCQ8Pbq4HUmTFP
6lmVOv/OVoxPjGLmbCrZl/igbGbhYhab7bIKzOMv096RtxkeG+QMVOisOAH9c6BGPUyJe2waA9+j
QsjTACC7tuz67zfsk3dLPzz74D1G7GNJ0UH6dEwptBhgjKL4jgPffpPcj5rrjTqFC2cu/j92NHzV
DA9PAV05ekQOaTrKTMlSaRUc8ofMITTvzfVhF7M2e7a2VZNzOhAQz9g+FlU5Lkm3mnrj70yWNimQ
u89vgc9GMKJ3sk1murZ2s6Ar7L3lAQva7ShNJbd5TEyBw+1HDNPa1+t1ZkKPnreJfi8AU8KsiaO/
ivU2vdL9X4H6DioU+TPgIKetYytaB/4KC4JQw1SIAU6C+fCV3ZxrIQb+B9VfcpLfLFBPg+YCnNSe
O7KtTLX0ayT0RYzaYTEnzmJIs6xvtIz/uhTPxxwjDEMGipMeSf6ZCnukOMnFSZzUW0VDQ+R+h0W9
3y9IkiHH6yjRiVH1+DJlxHN+5SiKEOm7xnNy4nC9DIIEYGk0nzFTeW6HyiqtKF3mwfmjhIk5tm3J
y/nHLfXX73S6ouxv3DVdgcAPr/y86UUAW5e7HshQJvvmg+nxC7ISlcH7Q885Bo/LZAb1fIVP+GeN
BFQs+2YHc/aOBNWXF+BveoG9Auu2heEgw+5Mj94GIBXSFNzOadc+y8PT8PzTeJ8huG1Wy5Yl0AzO
0UjFo1sG+dlQsYGikjbhczyBipLiYDvPYX9X1NYbj5z9Qcv5iINHUJU2ytFjMJ2PbgaOF6xybt7s
H9hjJSPbO0aRi7zM64hRcScxsh6O3kHrCM7VSjWB2mBd57U5CAeN8Z1MMRdU3o0rl8N6KlCzII9K
Wp9tgoAxf09BFAvU6NWvfm96Y6FUw0G4O8W/ukGT6iDdBVI+b4pURJv7CTcKQ7gwN9/SWDnFngWT
dcWCTQmhIh1YmUWQ/XCnMC7ksAuWIU5XiVJme8H4w53HMgk5URUTyH05Bq7NouqELopdGONhkFNC
g/byCABtrcIJT+BENA8U3cy3L34c/rfJbLumAMLfxAv7lln0E1ldrvTve9Q4ojsuChbRDM/5qSE7
AT0KcFk2NXK27tZSEl8fOlDhffB8886otSmpJ73zECN5+gKWrMEq0+Fwk2+ZyEq/x19Zikq6LrzC
r7xjwkTtVWP2xqUr2+sKehij7i840t1ilEsziNB0QaGXDSKol+/Tc6yN16Hb085ITYQ7ZCSDCq4o
ska1r7fuvnFTX4pBWW2N+BLUCTdtDGCyqI1/R0WUPPCG8dsOpu21DfDtKeFTBPKy1PQzragpbVHk
UbuDwLN/OX1y/VByJSbhM7eVmR5aZKxRnVOyb1DwX4zHLYjq6oqP47SEnx3befw2R/BnasOMU/nL
A2Uji7nqG4JBTg/fHQ2QzWPDXEPLARqwz9xmMgJyHugFiSid4yKuzCpNrERNe6SgtODN4UTPY1vv
iOIGEXhmcC3sQDirmZwobFhRho1/dBgxH1hXqWJuQp49BlAclkUGCoAknR0tTkkjS266NJJKU6Ug
AHoUXdRPa//iqMAf0V1RtmPWFNH715QUt0D10ZjXwBnlqhaiazKaXDGj6M2kY8QJmzdHIGs5eyoC
0RynmnIvJp+BrmffeqebjQjceJuhNgXzleGZVP5Axqwxq3QL9Lf4QgHyy0r3YCNsEmsdxhnbV3YZ
dRRaNbMkxL7NCvbMW3u98b7TWsCNh1Xzev2y/zkwpQYdrc5GY30H+RGtDZwRBBdvWHIWHeySfB8L
jG0CWukEC8NnDsWtaLeJrH/neevYFZ0TjGCKgdR+hAPZ6ZNo4Ff6GRV01wy+WsqT0u6y47QBMD21
oPiA7C1w/fTsTQTJ3HJpM34qKZUHHkIlAtl2rtBhThVFy46PUhTY61dCh3YD05x6Tez40tTnZ5hn
/vlKzeq6mhBxBYg7PrPN1WJL5dY6WevQB0PnLjGmmnrXk5W8r3KpfVtqODNjtLlMr+ySMmPztwj1
ZNZ9yBSF/zSJtoC6+3s70dDJoxRII/1pIcuAr95MwRZSYkq5bW2TDRWolUCz7bw0+p89WFiWO3kr
pjwwmpnGDitEgNGxomW7ASDoytLUWBR7CznO1IUponxs22A1ZUOKMF8QqwkVe6DjVC/EAmJxMznW
3Mre6lNjFHeBEtgigd+/SIlLyOdZemxa0OZ2CucN/Ueu0Ngcu8qv89j4QmVJt9MMVBipgSMUneE3
q2EqsC2ZandxGSHCJW3eeU1qluyCjNyUBeDggzH+wKxVMDcfgoa2yY7UYTzDf4/B1odO6XjApReR
dmghanInj3VOYo+GKmnBQrODkYUildNgEKdXPol7yD9FM7gEzzQKuO/7yzfXhY8oLdNS9SPniT1A
r7JMLst/10nnILBIdv1LfA0kZcKqpME/Pp/R/gZSEU42xhbyUp6n/dUt1fp/H3jXCaNUIC4Xw8ea
Qi3656pSq1yhLLrdDbjXldsevR/9kmy0Z44L/E44192BtykVCvaw9UwjwktYAiRaAcaoSgl+p8uG
E+mQDa5eprt9v+gKW40MtsRY50hMUFNV/scs02SEZ55IKTC+lHqucRdgpjasPTPgQrU8FbciM9bm
Pjp+TuUKWgPycwqtjjqORrWfDhg3dGS6KhiC3dVl7t222Mwv9KC2kcvrMlHlvCGlXduofGjAF0v5
meB+3SXHvVKDmiYsjGULq5RVbEKeEW3haZm7Mfbkj9zYighEr8wczrJXo0eJOyehDxn79WAozOyd
3eitRufYLeWaz6TUX2yBkIoapaOo3bTZOJkR97piC/WQMmIWVzcH9zbI2y0+R6du9D8kbxQBcJEp
WVrlNrE7oaAlpdaskLlr7I3wk3fe0dTEfNjF2M4KIB6zdJ3DHo4k8U0kvpm4oIitJb79c0jo/BLa
C7F1MyvgBFaSn3clpvOp6nRGw0bLuxn5zFofmK8vHZUALej91lDa0qgVcOZpGrXrNTpUcgKvS4O/
CC3UJI0i+1n/HrMwfXnUJLGwGx2FekmeUtBBhStF6e4yBu3UWjUmlhfOkr+D1k62IBR19HGhsPyU
SNy6Ki8FbnPFEW7Z+dsr3k5memBPfOYDq4GJUDlhjQLz1/WFenY4h82uy9f5evEHAifakguC8lDC
M69xm4SzzRx1OHAANz2AZ8IrqjkeAk1bdNNMl/ONWU2KPZ6kdwQCXGd0jd4lg3549oPAE+wPTI/U
t5DYV4lZfMs/UdIUslumOFp3O/kwcx10M6VbalTmqTwEY0UOubp6SqkSohLCaOYA349HRhLdmjBv
dkO3TriruBJceNYB5gvWwDUk2etHeaWH9+yT6SsYiBLYGO0LgHKhPRacSQv3whOuRwalYtQp7o2z
xj+6BaziHFzODezCwcFV4tEDrvPS8WU2AC7uHWjjaBwo/L+YvFsHJFpVBWN58Gbn0LR1FEoK/bPj
Dt7ycvcYlAM5YWbw/hVnz9JHFZij4YXISxI+hW1oInbb3HnErACUoy9M2vNrts+YwXSfEd0fKTDK
wL4Ee8bAvbzfBqxJrbgrjEFpZfJ9add/Fqk1tG0bd5B0Ssfd2B5fmay2ZGWBi6qgT67+e3Sip9wn
msYYfLP6eo62o21rqszGFuhxujDUl0g+pQ05Lfq8K+Q9X8VAA9n8Q+jCzdHpH2U2NohOCtkDpsK6
Dt3C7G31PWNgd45+dixLGWcr7s/hqLYFIdzGt/kPgyFZ5amPiGWfRUjakCMqLGn6KoaHh6msOEXa
uX1uCXPV8NlaNDygOEj0wrfoCgqTWWqnG/sgDpBIP7TLoPmkHVNyVzgmN+0kpH4FcsrFCGwegkfL
+FqscyTGGYTUb8EEH2hMYpn2CITDBWgl8/mKr69IZhRnXw3IDeH2iVFNoKkyug4qu0wTeS/SENXP
sW0mHDthK1LNydVSsFMORE9Go92kCJaENvOQdlbSu06t5Wjil5ySnZ1aw/EcVc0+1u5Xe1b4jLzX
my3Z3q2rOrCrfTUb08R/OpZUmYo75CtBVzr8/dkYtGexJ0yV+zdObZny66dWk/rO8oxP4SEhdx9t
aTnHtDQsazU7cWh5fZTOq9Gv/2R+W1gzJxmaqIAbfuhuEZldrRoSD4Y77SQqkHL4bT8h7OQrsEbt
YOtUaDNv2FF5E1tt21jGHfA/jyU0PqKX9YbFRhmV2Z6TJKmvbKTWGcJtNNmccib97gnlOY8TkBvJ
uwq42xTDX4wFmMTCOusabxoMax3mYZxUyb96Lc+lH9JPwM2XbDPVgX//3D/49xgUCUM8CK8aQV1Z
qHfQMIwAPUtB+tlaZFyuWteO8B6DGoSb7Ixg2kw4qdwcjsktVMtEU+rTnclSGdChPGB22VdUyoPf
EMgKEGJLgQiN9ojmbWGVG6eFYbscRSHAfaOeLV/Ei5cN+eT9uCg2lkCF5WC3WZiRkwCLh02Ogbqx
7AQpe9M77GxWzD80aYb3bChTqd+2bE6mLG0L+acEjMwlPhiQjypcF0poX8jFnnUqE6zn2YYWNEFB
oRqsRrHAnk+NSjcyxXLqlJSLfzx9v9gnvUO+m8Ta4YK868J0vqJ8291xrFQ7idGajDSS8b9K46k1
8bPrlI/VBVZjiuUJZ1+yltwkA4vDDNGiEIHIRF00DwH2Dsk1gH9NBYs44cfOYaowR0wXMTiHOJx9
S9Tqpjn0XLYy0mQpMWCPLOj5w+WYJJ6etn3/yyLcTlwluVs5p4MYy0Qn3YUjZK8Usvvlcj9qJC1u
/+rXw99jHBtwiyk2evVCkmpMwjE/M/RjwnYqjXhNMS0WvUdT+qaYRJZXgUueCSsRBH6VHCPyfD8C
O3umAjMTNobrvwGPW/sB1d6wF5lPPnWRReTEt3ohEGX/nML5zTnadP+1SFnOWVtkC0Ycc23cu9pw
yaehUPW+2mjl5r2qP6/OrBVvQY8o4wa6Xl3p9Mmif3LEB+Rr6cuQryeWgByjVkNESyRuHQnRfNXe
dB4zSw3NKb5c3z6vsGzsiFjT+ANFcG9Xh5UDiLFSdgcu6TMCYAOW7m89EIJhjah24SeU1hogy+eX
ltEcY34HLFhVJj/SM9Rj4dF0wBZ7GwUZ7OcXD+mN7BH4O3k1epbt7eKZb6F2zGhOyukjMC8NXsJe
KuRCyy1iMV2KuCfEZdXFvcSKzPlLQTEFWa2K7QtIyutB4mEfIqG5ePUyPt4wFH7zEHSym9KAdl2P
S1IZK5U29ly3IGFcgEuL3ZhdZhcN4ueeba6RuAeanKOzLgrO07IHMPHcEPjXSuKENc9UCoBNpaDY
DMBQq3Pj3f5CngO2agY9Dj0fVUSBhl3LCk2m6aLI2fyb2BXcUjkJuv4FaVTCrqq4hMBw8SwSm9V4
OaIv33qtSIJLD06hIE2ip8nV3vMyrbjOjBZOgLSxEQIu7MsU4NW4TJ/5TfkZp6fXmkCJXCPbrVMt
Q11TbcfzJdM+w7GD/8v9SK9HKpk8BzeMqwZi8P2uBTKlQQPIdlgv2YXyyksrFR8R+aOMRjo9DWyg
fM8DMXQe38ONB4IBp1w3dB/bfHpdiVitHvUIuwwQ8hAl9GOOMoALq4XYeNWF9qFzQ/td3DObyZpf
B2kpuQpPhU56lAaRpECe4UHWAvuo8nWcYpLOKibKjBotT++rcVrQa90vJ9CrrprcsRk4zODi7q3J
7OSIITAbsHr84gLUhOmxL3bnL5CWHWVs1pg5MOOOMSSpIRV+So1HFMAm9ZdyatX25BWceN8LWeGl
IJ6YMvXv8DlWG9KJ/JFkOwHT0S/89TaYeKlzCCNuZI7CuJTadTGri1/I5RaUR2Bfo6mB1rflzf0M
lt7hhevgU7X3PS/Rw66kt8+V0oCa+6zqqnf7UCimeFf7e5hQe4HBK8I449Iwoj/rXEMd8YEnCelB
OFLHJWN4gVQByDuhdwhCbPF9n32UVmi96cAJgXiDJ22eU867ABuk5ncUbFltZnf0sGF8u//LmDRF
cC8DTTUz6FQZrXTHuXicHArDbbYQRlW1gVkrYzTwsQTUGFeAT9PunrgDgCMTvgEfSUNNELEthsiL
uJ04CHgLnRSp07bZt+vF7m98gU6S8b+SsDlhaMZUvvdOoUHJcqmat83r9ROE+HZCuBAHMppY2Yl+
TJ3K7kqMkK8DflbnGMEwGV2OFFKFb6vCcotpth6RwS7aHzxr2WZT+GVsjEZ3IgkAsJTgKtXTb1h4
xgZgedY1hiOTj9FWF4ZItrM8UNBBlIaeeT+mHvcY5Y3G2yTfLPmEzAaeMoI1IsmYKlrShvKhVAcx
Mrq8kswHT++uzgVXO15YWQik6vsKBq75STziVDwg1gXXewCMmWuF+pAb++Ra/DSk+czoMpkyFE2g
ZLewxVt8dfaanm+7eAFe6hEe5FUmrJgjWKvrGKsJsqhfK0h1HHC/v2Ajgoff8eUDS9etpK0R6NSI
3L/SB3Hl908iKMmKGr8zIocC0DeAYi4WBFxsedxGZMRe9jo347Lad/VfQYvM42JUtEmr2kNekLb2
ue/maza9ZZIrzkMpVVOxn3Mf2Kt244u7auT0EsQHTdGjkHAMwIeFr/SBeodhMXE8DnVo8gtPm0EF
mvOgHWPwD7zcmqUYFqHahYdx5O0/a0kZQnp6xrKEnaIHO5NKAo+C1cYIutgAkK0sfQ/W5NwJYfh+
ZBVEwFM8FKnixM1bT9WP1ZiQKrOEPva7uVVtTFyJVIO3Tr6siiZ/9q8PFa08wg8nUDm3wbLWGVo3
dj2xb7ld/M2IVBYqo7i+G+FOqgCcf92l6lJy/c7gwF5dkZj8CjNlij21Vqt4I58q7p4qPK9xxGXC
uhc0myX2sUEaxvmTczCQQS302X3FpfFIv6nP3Vm/Ine0nsnwyakgYEXDyycaDH5battzoRWp/fQ3
rN9WrKoZPKtJlb0AXlON3+mIPA7TroIt9txR0+xQ7qa3+D+1Bikz24TV+Ph63ETbyxhB4GLng+xY
LstA9lucPumTtlSmCztuz6vr18dfznYw9VgghEmDXI1nyOv8PPqCNpEhkc0Rsxz6ktTPf6fJBXNE
uLPUNwn1FPBQe3PGJeL+Q3R+2X+111T4N7eyWJFRpETha7NWi8LOGeUREq5F16OQxak78LdBQzDA
Bx1OSXlTSpb7JQkkePDeywZ1g90nvIbcASQL7kE2A6rBIWVquHiXX07cZDiCV2OqkRyRaXQNRIAd
o0dzSrcCJqFMf5+eJ87y826USQmZQ8xWGyjWgTqqptI/FGsaTtJHgaaOePv/AcVAuAd5QLGW2f/p
GciY1gh3R+CLkI5re+6WpFjnVDc6Urzz4ZS81fCwk3JSTe20CQGJBIszuYem02pPhySAqDLmWFvQ
hNDPFKqOeDrkrOMFoKnd7ZcltIJtrfq+SMjVxyYMmfOe9VWEKE/oN0bRXvyVUVZYzUEX7UgnXumo
WVc6r7JLIauNt3pRU9PgMP16CXKjqcGm/zePCq2bODz9k7oC0mdlo1bIECWwFywlNfaBfSzM0YVR
kMJ+PXqKNu4OdEH3/WrGGd7F9paLI7ZqTgiLxWDcRa126waPOy70xeOXyV1CjTL9VY7k2BSHSPeC
HX7ZJhsDWqJgmyVxryrWOx1WZwH916mGG84hujJ3cpFCMgs2qD1J3R55HYL8wTXwDnHxr/F1batk
cf+u5z7HI9WJNI3kobI+KEiNFtfoBZQ51gqyvFFrX9wKtKNyYX6kFc9RhfqQsyf5nn+TgjtZx6Gf
pdaLSB+PwEZxHRZwbHZp9iMIrokRB3gjo3IRpPMCYzzhCln76xWNNYLmambEz+Fec88Z2bRV1wi2
iGJUsvTqHU3pdP9k16/QzX/o0FSa9wkbsRFMB5RpDe+Iu0qQj1TAgs7Cf+DWgILipBCrKoyvAAqI
+dMQxHuqGGGXMQTOkXLypfkoC5jVhFF6OSk7SSXfPE7yWSarJysXLBQIjDhmb6OPOm5l1Eg6hEof
zshAqpc2IpJP0MpNl4Ux2AKvfvWvVZ2TgGs3uURrJwa9d4pgGPLNpPUNOzcRqyjff/Gb5hNEAPyg
xbYgaN72TNxKhqxK2rdJwQZGFidHMZIbAGFXF/2GGY/eUw1ig+can1Hl47+3reo8FFAslx8hl0vv
UdmSTv822Ok69ZtoB/OEGwM0H3hZ0mXbZFJC0q78jB6Ko8hxcT3XeJ9IEiYbc+e87j6FAwCiDpwL
6jvZQjPR14wp+lyzcUBVdt/NtBk1shJeWDb8ytTqxEPTGRIjvMTziVnudlxacr1CBt1YISs3etim
uh4kY+h4p3oCXi6ZzqBcotQpGTBGI/nW69SWQNB/tkOwrGo3TcpN+794YmLgsxEiNM/axBukS9Cn
yQbv5eKlgVAw2B5qHv95yCdv6mUsyqgJYplfxcbs6wE2AiFSe0paARgOCKwABSaqSf7EUgqJgAS6
VLFx0v4905iHqmxJVroa7smfyu5FErh6bgCcKdUgqwGj11cR6iU96dtJEPPCgkgAiVQx4IKHHVtH
RvABItTFje5TclVECosi3yTR+70c5o4sm5uMMRa+jQj801zjB0YAqSX3s87DJ4BqOtSzT3wUwmQB
US4/1lN1p8uMzlaYYETrpf5y1+TgvPqdttJgOQY0A5ETy7lgnKsBek7ZySF2lCBkkSo3ipzKR9Lk
wEvzRBfo4EaXseT3rIzccFDtI3KqxZAdNo2RV7wO/nJjE/JLREo/TNRJFfnpOZACtj2Enksr9BXm
pGli2H27bF1eMFUkLxFNZQKijk0XQA2ugUnGhhuJx5OlY3dPF8MaQdy7bO3JDEL+17sMPuMME6tY
dmx3eGpML8sWlKpjinQYNTiJpzJfdsc/Z0dkk2Igcu/b/vJW1TQu3oCZ5iIdM6zCFX3sKAOoWrsq
dIBn41PbKNylIzCABNEhlgjhb/mR5AlClYw2tKEdW/ONppkPDiBHKFEDq29M2LS+0BMyDYKTdIjq
UQ6E57n5LheJqhBaEDBps4sLoR1kQPUKsa/IsUIilWiHLCyPhKYv7AHhk8oNVQrX//nv9tsNrCC0
TZ4Mjb1EySvY+5qKLRVjZqFiYrYTsIGJUcbKjDATQ9zq4TM55j+15ohz8S7PTaXlMYiN8sVSkB9V
Nd7bcawiZ26sYybJX7bgjiRn4K4+4l6SbSM0FpYXje7uOGT/J+gDvJKgBrzve+e9g2N7tk7Qts+m
snWBk/j0BqO3oZkuSKr57nvaEgfccpVoFPjRpAUQG5YnnOS2ROvLk1H7LjOA4j2jsFwSFghk3wx9
xt8KLLhYKBZcHDIQr6Em9hIp6A6QdgervLB1/WC1dpyOIRxf8LUkfEdiVk7u2F/nwfbOei5PMcky
fb/si+RuDh5P/RqoDdQT3CJo3/2OyIF3KOQWfIzATDREOXcASUV9r2cAAjw/Q9AMmDz5EQCiijW1
6zTU3sAwOd2UPXmvt+E9CJmyNzFAmCkMRPou9EmzoGqRpXKLC8SAP1cCkFV/wKwoqbvoIaJUwdYG
0ROgpP0MhyrC7q578wWMCZCJNkjbjyzGCZCBN+lKf5MvByglttck037pKOAuooiLm8K+prQfFLQ8
mujVmxJjzDJqjrejAWtXXrk2EwiTOptTKEdznXf+LeHChTpBPCGDQ2Er8Q+OQB6YyFvnC8qtUlJ8
obFM1jp0LI3+Je0HD+ZI8KOJQHmRQtvgM1HQJaEU4SgH1IsM9WjYITHbOLFUVZTcyzJoWVIxM4dS
TF6gU71GzZE3WdMrFjfi0FDX3bhmN15M71Mh5kIfzSWZTS2YNSIDl00hwMn71X+0CasCvLnWOmTX
NHjxtPv18PwUN+Xk3s0FoucgR4RBjq2325Ns1GoFKpIfBxor5RM6osiTkWVqhoYeqmKlXgaBhvSg
RC1CM4Qbhc639ZuT2DR11uKFjDuUXx2/DXL23IJb+W/pk8qHEHdPZCC+WaUqsNIVG/KEeRITEbcv
Uuhrz2FAwkXNCSMASvcSdjGouB6kWV8cuOtRLZK/tgmkoNYj1WR22doQOG4+p7Kkj8xkmWODChv9
jkJWczUCaRJYZoVxnDvS0Glm6bfo/V2qgSBGYZGOd1QX/AME2tNtQ7B6jJ0XimgR0DR4/EBrQgB8
V77a4zE4nOgklYxHxmKDcmVESVGf2TxuqqaES+zq0ov2itE2FRi7I++MJ9lSWuXVILFun4A6q81s
iz0zlIpMrk4Zwcv3uoUqR/FSSGL5L4yb0Bi3IEF38m0muFuenlJb8zPhW6FVqROBW2WOXrvZJ8iW
YqWLPmJnEWoPnLSPm5JO9ToDm+x5M33nRxCtcfzardj55yCfyeP6tH6PQ96Kl2DUuyLmoIy/5lht
NTUsZlbq9Ph3hnnUbE59C31HCaUEj/wBuVpjbx7tnkzzA7C8+WFqgg7EL9LzhcSsm3MKih/HvMfa
wQmI7XCB6Ax/LizWHMZ15vwKg5KI3/y+rtKhxNNfyP0dlvOgwI8BF0Uoipb7XV5inzy7sA2qffOT
+daBumNZCwZ2BwxdaNUk/aBqlctKS85E5iX7uf3fC78LBIlYCsvaKdeOJz4l4gqfq2SUB5L9R1Zt
CEm+puhi1hTGB7/Do2l2pjxnP8uLa2yWJsAC4U2fW21YY26GkRGT3GUZh01GKeZLKfZYPFsSLqXH
Y9RQkPHaWmU6X0VL1zlcbD9xc+FMqkUdPaHTJrntc7tIR/87Syj/10p9aQ1CDOJzXiO+XMRRh/uT
DHJzyk+u2d0A/J+Mevl2SXnzmAJ2c1yt9P57QtqnfxOFpFA7mDSEZ+tPc2CicmMKatPlRePzqAfD
nHPYHypbziX1NaTd/b3REcC5V/EC+V0V+3PObTYa26x+euOrxAGF9sOaA2ylG9DttF6l8Qqs6mhB
G0GCQEODcM+2jo5ulBeA7HkoZc9jf60W1f1Tna8EUNt+2z+FcZdYhvyoSGBb7M7iJnaDVO6EQn9G
ddQmmnJfemj4Bnxxn41EjOesbSpqM9MTBQtzDvWwirX1/0+hqPzio4cIgkxwPwqaCedTqXGH/K4s
W7rgWpLuSc03BCTVkL0hj5wyTFbm+WR3KxVY4xDG9ShWSPG00FVhyHVrMkhx+HNOqU3h295y4Sxx
DLkOTsouzb6yzMfs2RTCkD8EcXVRQ0IEwVLZnnRvcGdF9tiF1vpwa8+JEXMCjV0dunsdfC3SrBxY
n3xzdSESrpvCyfOkW8whbpPAemONa7EhzRuKsTI34JApsyUVIkTu+6Y0kLAAc8sW53XBESWJS2px
GxmyIqlq3+ORbHcIOM/cnnMVsJqrzr9Zh5AHmOEqABVPPqI0g8u8msFOiDBiVBGQm8UhmTzvuWXt
7pcMy7tktLWXLtzjlKlFwdtikCE0dDBRyG6rmHBrSebQLjptbovo2TrKXzqTflJwpMc49ir+stDQ
Hqhg82aE44hoCvXVZYddYx+4JFYH+SH089f1iDLFrLsGYdwDuJ6zYDqQnslrZqNr3sPqkJHSZdL4
P3aeO10kv7pmCzXSlt0yKdcOAVlKf473NBGuyL1p6DJxXQV5ZaoFkM2Df/qAWSTIwbwZRhYOpzTS
eRgwZ2YQJKgvzOHWpDJRfymOOulsSeFdw8phkV8n8P99Ru6QO5t0l5ZzXgFgRvKpH4hVHhXNlXpl
0MnmHvGa3k8bXLI6+UZ1kRxvgFYDwjtdrCR2XFDAAzX166HFCWFUesnAYCGUtC6cSF+ECA2ZE6YD
JXzfvLZB4vu3fbzrQ55YZUuovFgCYqQAOqOKHMij7AaqjWc4ajJFXRrU7fYFbubNACijNvoPvkaG
IrtpIPEl59roK+EYyTNJmRH+pPXn0vlLcgVNMRwKOzNngGxOJw/mK8uY1ACOT+rKbxzGdJARJBrD
3Pj6lePpoBewjhW1O8MkesyRbqytWSOZmCuvGrRz+ifORabJ8Q8kdo+Kd6qBqRKM/7Y8FMFWpeXj
VwOX53MQh7gfFbbkIHPmE+5ZufqUZ+Tf77SpiMKwsznxv2a/acT2nan48Q+tumbHHTUdjqNBhkHL
gfaG+5KKtf6k3uMmaE9Jgz5FPNyEefoJH17b7JT3IV8r2kSwGOiWReGr57E5FJq2aakqnX2VGVuy
OhpLV8Xg6q46vafznNm1l7ucMq9ZTTZvUJccQrv3lmmOd0tUWbt5p/9zsg0GoIE9kfHb74f8jJ2B
3ppsGKib54k9yCCbOt3IURGD1uObJ6YkR0DoK0uxUnESR3Y4vDRAkdeWu8aZr2xJVh7MTSIuUXm3
LRhkV4LI5PdE6SYdbsSOB6YA+yGD5Qo8en67mhsoemylPrIV3SmNBUH/FwsyBSqqCOPliE8CrlNP
HxPMowz7yqN9YWI+C5YwIPrBDZB25yKEfbD+tyNwRgH/ZsTOR+iQxEBQMEE8p3HpEXQAYn684/Er
90vqh5U5hei+n76wNNxhShYmexVKBiNyuTRpDakVLnqAS6mMekK8xf+Kkyras2J/yjUPjyI49mdb
RW8e7Tg6A4gwZWT8tPbJZbQmqcWSfQHWAetbAIGX8jL1L1AqcPTlXbFk6ImiedH2cQngCzZY62AQ
MrmxJJbEmVZ/s37tFp7QrWlv+fsp5lDq9RyWXMRnjSSAbGUGeUP3bzl4YHRsge+Pmj/noz/9LbJm
LjgJYYskEbwZWRA6Lss/iVcRo4vwCamF4jc2BHMKfe1izfFnULBeLQhlRFYo/TTJ1p3k65baAwvi
2zdyu5zmuvIEnzwow2BR+IPmbg94JEfo0siNc9EEArpmfkm4nX+XOime+KeKTXlBAb8kpLyiWss6
eezL24DRwwqoLD0GGupplOS2rqcryqZkyPk0sD03BZQRxadDdF5MZL+AZC4RMkKjn7ojVHMlnyaD
gILNVK74D3nq8HuKpdB/nAG8AJgII/PdQdxWrwLAf7mOjjuQp715M14Wc14T5HtVnaDxVc58u5a+
InAevcxuAaun0JJ/OPI9OIpDCqAiZQ88E9CG3p6XhkqwUS1mIprB1xIO09780OszWU9JPeZ1itpp
tXsjuWpQtDXcV69DKEtjq0PLHmT+RPA4G1Iq5P67Gh9F8fSSAyYN8Bmrh0WIM0plmgIZyOr08Ifj
4eMsTC74Q1uy9Iuq3rDzyFtNb80H+eG58fjTB9wrmw6FSHZQBtABgWEhVKpBoEOIiaVnzrIELSxk
gk9FKI18Qma6TRXdmbjYmZ+heFgqvbCa5LdriaYIU2oSYlcGkKz+Ol2uPz2QcDNcsdJoNlH6zItu
OX3hTy8rG3j0w91p1D6WZO4sYzHsR6+Eg3vLh2gFmZbxs1mcLs12PFTz/2NamFAk7/0l6M8xWDvz
YoT+n38gDhb8aSwD7qOF29+0D7VX8dkxPQpcScfNXsqjp9cOkuuuqTLoFreF38vaOtx6z6gUjurv
L8mCZII7NOt7++Hm+mq58+qGBtFF3cmom22gIiLzmt9P1HcTvT3lgIHVmU7vgglbJLTcm3p3Q03K
qWQOX91MgfF0HQEFAknQP4sVcr6xCOyxEQELpeaWy3QN9rzB7vpNcBVdNdtNIHPzNxjVNlJpRrTw
acyvQrJGHtANOm//3POPERhq+0GcMwXFU0161xgSJZxn4fG78pEO+rL4atZ0AYs3SF6/jWZtK9TQ
nlRL66rz5lBvFUECx6oJ0+iVvopf03xjOt6GTM4Us8j7bmk4HB3lIcm0dfvYM9ha
`pragma protect end_protected
