`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
TiYK4C15B8piYlGIa7DJss7Ef7t+FFCWKVkMYBCbD8UNWl+BekSBnoBfgKBlx6VoBRSQ0ltv+Fhq
i7Uov0nYog==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
GESg0XHM07TqdC2ez1+VTv8PnpSzW0vJmnNE/3ZPyS3PY3eWSKhllEib4jkh2hbs4xEebEs2xbDv
iEvGfd2LgMq3QuEcL6ehSFovPqDYmUZEsA1IxvzZzdJoS/Tl43j3R9JxAYZ8u0OlTetp2NINGyOw
zwgRLLEhdiAC/tXL7wM=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TYkMIORM1zvszFJuhrcwMNyYLroVI9uKKQrXJR8IdxiqsI15b+q2In5U1nko7NltlSKyz7zaBkQd
jCf+xXdlIzqkBGwscB2rygFdaQWku2XX4EkcpskpJWZWlrmE8xfZgiKlCF+quFgf6U7WPT6QDSuT
c5vCXsX50syC+73qwBF0tXvl5Kekp/3ImtH7u8vufi57ViQNfsm5F00PtRw+Mkh5KBTFBdJp4fmy
4pCyn8reHaLSQIezs5I/hVFr39p/LLTDjjSDTxmbrGlH7TnWwq6dIeoZHr2wbfRUKbWGPv787AOH
yaQZ8Wx3TM5Q6kRIH0DZMVIH+E3MedpZoGTfkA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
rCWNXSw5sBArI8CCDWVtV7T8Ng7ZOzoAw/Y7Xun9wwH6oIaNNKNBm0MrV8tayEoCsceAt0GUssPi
4qY5kO4FSjLzhx1bo+a7f4tm0ReSt0N9DpB1q66qg7kngNaeX6hIVhpKENEUwKQAgIEAG5xWTq1f
N2wUw/T6DvHUvCVDqYdm2pTQ7u5WfqQ1d3iNT8Ga8kSbLIecxu4nX/j7DQD6R7Mlp5ZdulK7FPOY
Pw3aMRDFDnnHRnpz5TbgIlJ5fns4VBx/76NeJclz2qZNvIswlXMKKxr8+cLnHwt3pfKijlA2sKU+
T+MB/Jl1/mInXVez2SBBn1hOpJuvEnSbMfKuig==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
c7I2s0FG6x7SOpxCOzkj/nm69ulO13cb2BV4MxjYNWuGj8/I5Blxr+SkfjttL8OQI2l9mxAwf918
OMQB4mMs/Rc096NtISZY/X2ZGFqsyJ+nlm2cN3p/Ta05u1A55E+0ohh7NmyqcmStgHfqpOeBSZJr
0/ll0OI6T3FqPvzw34QIowlYHotZScvVNwDHWW3opqhKeaCNhBKxu2S6Ihfm4vTvZWHYQdeikpYm
qWgrn6zQc22w+HoN9AMf7X1ebLQTmUtvs7wh0wCaZJ742pfup3rJEEidr/Rvi6RXFJltikm975DO
pOIdoKnM5Y7Ymwi0Tj060TcmYPMwV98Jh6GqQw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
CtJgYj7Vb4aQmN5ggOszC6GwUJr+BDcACzcVkgMbUilsioMCNHXHudqWUtMsUcQtjhOWMbONZw3v
F1WMSGhDHLLNC8klRVrZvqNyPIoJPBTFrizzgo+Fbxpzah6AAE/RZl0lkhtKpGEz9XwARLOoujkT
ziopXrZz5dXYDtz9X3E=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
DMUO44MhwVFFJ0AJZpYPfKjkzFD4X6Mn3N7Ymfj5c/Dr4mrE6w/Pfj1L9WebkcAxBL2a4gU7SVjW
3izO1jPlgmqP5RuXkvqaN1gzwkx7pyQwyITc7/kZZ+DKIOyRrpHLYfUSD8VYmIq+abCwgS4VirUP
8goYWu6DZA9iO3cGMrlM4xQ23Gu7KyP/SfmWfT1FeS1XiqV8QKC04ydkUpnUwXl3HR6v92rWEFiZ
bXnUTICCtmgwZRzC+04MzZH3/xtsVJggm7Fa4VT3hxASt9hvLpb9pdwd1aIZf5TKJf6W3LDtmG3k
LVlFcLZ0sjh76CubiukzzF1FDzxFET9BB9NQWg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 151824)
`pragma protect data_block
BEbVrHROuvUbO/Kg68+QjzvTBAWyi697rsX6/IPm4x2hlJJzj4Al9aIZHkibSkGoRCDAOI40KHrb
VvqE1Z3NpUCuOgato7ukKF+q3N/EEZ9IiJk7DUTBE+oNIexjyde1hUHrnKAO3roVugTWBYf3dB+3
3e/97wZ9oG0GjiSvwZjss0jD9kCo7+5qZNniVrZexHqLi3dWVPkFt+Ykd6PBznhXeK0j4Da6ZyPh
zGAypv/6tXS8vgwm9XJC8p/AEaD34lUH+VG0MlfcH94kAPO1mZPiHf4SnRO0y3DkJ764tdFnMDJf
s0qCYKcuMbV93U7oQqX8U678mc1fY3eENorvlG+Lf7/IPW7jXZrTk0LwyugmLgWkfREw7IpVkJtC
w4Cc2lrJ0ZWw0mS3IrGBX6epa4qW7YkfS5lSKIWf5Bs0/FjLGkAu84oBLHADG3qRNQdFGvi1+cti
yNQ3wT34xoDWknCafd/hRFhkKJ5Fmr+sC21Q7YtYPW1f82QtfedQ54zrPe9F3mA9fOGdBSpmRkMw
mveWnw72Z0a6mvQn31l1IX15Pi0uLUu4kHlnbXB82s9CLyJuftnSdUsz9GLpcSoOzi2uuWCgsovy
I6AcaUx9kOvVi6lNJqCXpJQgTDQDXySdKyXkoF5y5daJx7LijxwlZeGOx2Eq43VXm2RImyeekdh3
Mx4mCTsdNLW1UAS6j9qwTAttAFwdA6qOs4GKGvptRUUk85O0NQDFAYsUuEUD64M29llh7oS97+7J
Zmfgu7xwv48kRqJ8JZxqivoOTNk4EjDZD8kEsZogYPlF2X4nt2pbrGL7n7lt8nDTjvyNKP8n55g/
3ohfiDq3Z3m//Qh1nulii6wJRKz+wb8i2EYgR6cgyWFmWcfyeXSH0cOIYVdJR/jFb9qQNKeZXHM5
zjbCTd2r8bhE63dasV5XAuFW8sSHltHtVW//gVDrK+cFwdDeXoiTygH30nXSgPWnqAhNXOrGiY51
P26uGolMAkOu7Z5xLSRCTaMbw0sv02Ebnj6K2G+Co7KNAiqcEYAuTnID3DkCYbassnsi4jnSoYz3
6QyKYzsXhg0lVpZU7XtxtPD5b1UzChssuIeJLiVARDOZzTFsT53kySQwAG71rcW1VfJABaHyJEpB
FR+wWiQNrUzg5aoFDFd3ilVVG1nyRA7Y6r6S7Qd45r5YIGNXVI7SDXX9APiw6v3ILkiHyjxJWfYL
A36h64TUOkj2bAAGP8KBTlARZkBPfTXza05PZBTjZq9hcf3sutp6zgMWVYvUfb8AA4No34CSEWYK
wIefkaHarECLSxxPK0iMnYlAHNUX3HV1JfNW5yb9bmFiE9PLWiJcgOBYbPnCzOEn2WocgIjIe7lx
HOP+JviEahU2aGExhSSyHC8sQs/sg2Zg3TWySx6MD8G5h6PVujT2fSG1BsGBDwyuMHcXTDCAbzRd
KssLLLqL6oMPpn3rbdwKWEzePCKISHks3RGK6nYtHhv/JxMh8opmV7LuelEH1aO7AgUQ7CthJhL8
qZZwP2Voilw1g6xa+2328DzZgekiC35dEnkP7YFN3cBturB9S/t9G9lw0+8djBH8N9b8gf+Y1+c6
5rcpxeEs8q7b8dKKx295SKCfZaNFaO2RKAwfAzL0RjkplZsrdlHYnJz3iRRd5QmUKA9ASgmDMkB9
ehcYUMzq4XrRc+bonZZmOyproAeQGnRAaDLRhnISuK7R/bcy85m6n12G0lZsDjUkL106qXQreg9j
xyQ5sSpX9G/JKcx7KP5GEw2XD8oGIuVnOjPwZUnigkM7TDzVAsJMSp/F8gNWlPaH6usQwgvHu4Pm
lw43fFm2wyr7/uFPospaWdwaz3zd2Nk8f2L04bfzrwGb1bXgl3AXiHLNUttQAYFnf+Dano65lc44
HSB8Lf60W12A9kUxwxYk1Hes8M9QsX3l8UH86bFUwlsF8XgNrLsrjPecyWELfAnXiRGe38P1LGTt
3GJakvaKTYhkq9HQDZT3N1RSFqwpRpZGECuadwXZcHTubv9BuMliIQv4aMn0xM0Q3WcsR9ru77hP
F2tPNqE6YlSDvk/84MOJwgsdaqR5tQHW6ErlTjb1z1IMFHGx+rtfSdVb/HrgN/Bnpr35gxM0xXsT
Wj2yCMBfylFll1Ix8iLFxWax+qGOWFlDYwEXAD5KWMQ9BZjbB7QZ5mxTd0h3KL8mjK8eOD5gipNc
+f0DL2jZe23Dl65LaAe05/+/r8nhw1bRlZ2r8hASeX1wG69UYAOi24L+GEprM5VBKOHcOXo/+fOU
vcUp90LNnBtnThkWlW58D58pxox3B9YYNhhZ27716Kl4bPc0wydePfVy7dXl2wRVzosP+nnmcLY7
W5nc30GGvbQP8VnyWPB4S/C+3anSb8FQcwPenB7HFN9DuJO+23njFibL39Swt7Ev2Mqlsqj9Yiry
tDXMQYSlNWhJHBQraESaBrz6qJFMpC45Y/m6gL9e+v8KrCet5RgoH+cVpXkInd/2fYD77kZrGVfd
QrEnS8SGaAcK3DcRteMXoKgJR9P8FasCgMB26sPqboSAlKK3rPYoFns2UA0fIii4GrCL9uB2pi2x
9m7RRk9MOOaHqex1wGst+pbfy922ryMp8WVnw0OjWHUtxhdPt0LfVCtTBDgj2BvVWimpdDDHI2O3
KgBEIubQYOI5VO+CI4H6HGIWHUb/sg4mqsKwkIWxAwC8RvlxuEbltrnwWK2DLAsdjh4iSGPCFEv+
N5LMj/iGULSw9h32t9VyGh1YAXMB3On1Opay9eIXn1VOgQ7YQQDK/76gPIvy3Icz+7wxMRk3T2oJ
3LuUEUyCXXRs/ahwZYhlubvDzbulKiNOut/VpmEovoAP+TNsZENTQXXBoye87fccV0rI0gnqV+dS
HIE+YV5LX7seAicwy5IkiS+ij5qYFGJ+O+mccm9yvNPkeIZ6nNB2xsUJv9Zy7TzpRED8VDjPF4ME
EuNAApGKY1Zguy/BD5s6O1M/EgPyOkAdYMJVqz31bk9gdcpjl9iZGeVolmsfiGo0sCUKEBxpDXXI
ZbNnXoJYRSns4EDtnWuQYGqTxkbZvw5Geokf8HqnTmksOWTN/msHN9iBUQ1wv44fCKwk3Iv9rn0n
XDfwF8yakvJJp01qVs48DF2NeE26y+r3KusMVJi59XXN4WQpqVXWh78aayqKSeJEKHEbs/YI2tr6
QeT/JFZfYA3ct4jP0E7A4tg2Ovdd+54qYr92Rjcy5Dgo4jVrNSgO7X0+5cpZAWfAZLLcl+1Vi4Sy
hfxsJD1DUfnDh3Az7D1CghaE5bTd2IbBvRphHLIOaKCnKYMiUw6d2Q+bH81D2DOlEIptEwuyDe/T
/aJ55xpLzfbeiYq4yAKq+p41p4+sKAvhVu0PSkODV5O9DqjbLleQyu31Ue6V13vbBkLyCVdDwGkW
YHucfCfyL8TBqiTFuwIVK498WDfrWg1rLpvVIZceEV4NXrrRRhNY3TvQz4V36S4juHpBL1ddXO4V
r4gXspF9+VdJy6PkwF9XSWv87g/EruB2lSY8JC+WlgprD+3cmde5j8V6VKc79uHPJ05wSzSITKSg
thv1+H8Mwap3As3aOdzdoCqAZPO8K3iLnpoAJF7frtqo+FXcsFDLZu64qSFZVEjx7L4HnC3e6KQi
sddjYI37oQQb7++N1UeVl0n/bz4W3J9TOaixG6HUouz9ktqlYc7KuyoOOAFNgMDRU0AGOfAD6er3
MW1b8ZsRxrTrXrWCKX/9pLjqvSIFfj0LY7xIAaO1Iv9eAz4KCDHHXqM0q4k01ie6CXtDgv8xMdLA
eX2olDMDmeqYnRVXRk3XQ0CLNbypwkbe8JTzag7K085pBLOpzqawx0uIGXSHwVwUgneyy97wLGc7
VdV1cgHmeJbZAUIm5tA3hwPEVksu6tRIG3VXnt2u9SUIJZiA/xAoSyEpJ82Vrt9GTNoLf/HVSAkX
tZ715kxNU/w2w3j3cQCeITln0zDSObqwo2vApzKyigGsBiGmLAl8w277hYHcJa4nNR2UIW7Ojvy+
yJUlaIZoE1xIyvfv2umQn3zNLvUCvSuCeY8V70I0OXT6QG+L3sBb7aBxTY9upTCsLh/sYEbz0JPR
Hqmmz9ymqRee6vb7V4rHaYwE8rWCAUA7Rngxoy3TxbeAZ4R48+ovz/BL/pnsH2aSq+MTVH2vY/BP
4u32HXkSTUcy5yeKUKqukKzSPuI0p1xb/09nbnwvAsuIZxgbb6kog7xlZE98xFiFHVF1tv2CCoDz
gAAK0J+CjZI2wkPPec4wQQyjTwnLiAbPv+S+xuwjDHoqNLnjUyfeS+qHht44w9L3blAMMoVgYfGd
NO11GZzyqbwChACQEKb8ri0Pg3isoQc7WR7uBf018kvjKw8RV39j4e3guCRO3s1FLgwUUv0Clw7y
MxSdfd/eqTKMN783K58OZxBKVOyOgyQWXgq73Z51is5kLdpvn5MqfCQ19V7ySNbjeMjLcyjWNrh5
1o5Ly7/Idqks/pxEtx2q2oUYdFJ+QBLIljkSvUiGs1RfT6MG86kWiR7KhwIupGLkgAoeIIDIkwvg
E/Z2EcjfqlJOoA3HdYPfe0NMtGvgKHyeCFDNK1eTdT9QDveKUj9oZSBRg+VpuA16pLl3lsMUzPHM
b2DotMpXY6MRMWsFM8hrCJQ7jSi1koomjKk1K4MudajzobHYISi/ucY4wbhcXPjy2wrYIF7+oVt9
UEHoUqGTxEB+9QpIORel3ne1NwIGJBpOr0sR/6fIMjspIq7Pq7wYn4vcneNNhUJbW+YEzqahnNZY
ad1+QAGREXAldYe4Cw2ZMxAzdArSmHdo7bVJ7DHNEVwK/JmkmvtrnxSHwNskl6jV5Uyh8eNuI9r4
iIqCakT82ymxOmDtzrI3klnR5GV0d2bKB17tzJol1DIkZR0eeeQSzLSnAfVd6pJ2lBwgVB+7Mv9k
YnieRETBd7437GY7huSz3xPBM75gnVwrYhgsIl+NAuzwgXOJGM4p5SJxZHST0o9RZ7ZmORdAdGdt
5OSO4CCcbgG6cf49XSLrXblQ0uGUcQkrQFbX7MpkwJ7vdvWV0jTSzdHWPacZglHYEiSZ+Qv9IQxC
PXuiKXjpMzmYZiULrD56mkCfQdJNG1M1FIBqOOFkQ24/wv/FjURFlXTnvAmJzZKzMyKH+2gH7dZA
3Tf5wjhZy6oLO/gxr10UAnC47VZrfaXQNLUegmuynpLQ0kyqa4nKWIMtT7gqf8TlXz9UbX8eqqB/
wm3FOX0g9sOKDUz3/iPjwSbwGuMJu/q4i81plZXIjevSDQ4e5roHcmrPwM5RzupGPb46N9lHai3g
Ov2R9jV8RgqZLfyQFim8CdpwW3fIwaBVbzzXwdj6idxwrVh7iJv96oVueoIomzC/pK+a/ZzzxKtB
0yBHP5QqVGbFEgt/ts2KQGmKILxuDVq73pe+FWveTr1trmhCVlzH6tH9oNLbSMA47B0N6ySe+nS4
wA5RNDG/sa+2Z8mzIKRRfdGq1OqMyp4XHYr17Yk2mXUDVCII+aglYMq8ldUrCc04OdDleiRlaJ/G
8Jml957V+FYOSROp7A4qs9CKbwbkQ7FZ9I+8kTKa6J1NeCL4sA6V10WuRVOnW6DiybLIM3r87kTL
tcCLttrB+POOG4OIYnepurUshGA+DNAs3jmxFSZVzAd3xAMwMLXMilV2obCKB15b8frHmRoD5L0w
ZH75yGuy51wsQGtiQFpm3RDAkOXHl/Lzpd+wscBD5jJlb7kEWCw/r9bdIVZ2m2m9QIXOh05dN+dj
/GyvMah54QAo1mDe8OKYEx78JgKqvspCso97zqSK4X8miErY53AEEC1pb9on1icqBlgk9ME3DmUm
xKTBzefm4dOOt3FrHJONw8v59+4alL9/DCaH7RxQO0YG2CN2MvsSS5PGSk4EaDRS64WZMS3sD7fj
orHRQWxh3YtxXBg5uCS8BFEd8nknv8CcjuUhDJU8ZbL0BOwKx9BcZ/uJcKxZHxlMx956XoL39twS
r19wTOtREI4FRRReFThwtzwKGNA4Bif8pLW+fxL5ka2mak4/jIINTRP0OKLN81ILAVmyKxYtxeaE
rQhOwMn6o3zo3DKAr0I60JyyNrz3aDPOJyVe6N10ZeNNhyBHuWLvcrE2/nIlhmoN9EhdTq1wlCTF
GyNaepBpBYOeO0ugnCJNQ1NIgGlp1BdpqZ1idKkMMS780SVLWDJSV5IKZLC1SYVdM8VxuccxyCeT
wSsqz2xzsQK2LrWNQ2BZ6JALsCGyEiVq33cJrgfoegk1qAfts/DR/OfuAuB08W6hlCaS2HuBQi4z
xbYucFxqQ6BvnK9qeq2jvG4dDaUkRYtcNev/Z2U7k+329wPYzbkMgyXNAhBO5QVzX95uy6ER6/sR
HpRDv8cVPkc0yHpOlB40E1pytfRHkip9028R8EXD4yzWVYKcuwXL2CftOmFcLe9at1nVv6CxxvzP
syk7G+sk0lkZQTJOIjJYaFutIXuM8KRoovO/Se+CqqxAmtqJX0QqbdEZ2R4lR9f2Hj8CB8RzjVyP
ROVgTNHzPHBjbEEM5ipqK2hT9YwYiRs00i2Yy3YSDXBtytbIoTmrDawNL3m9cZIdmtN4YwUAGJxT
9wrgo1OZYydgmJzex3hIjTdeyJiHe1HDLphQnLXsLFsYoHdCfUP+JkrXsM0efEJk8J3n2KDzR4yN
E9fcEz8DNW52pW4tLvNpE4ehRjO8KV5yyWQp3b6U0erEudsWcmLcnsqZ9QlppBKArOtrg5WwUI3F
FeBepa1ul3jBEaUZj/E5Wfy0Eqxuwz2PBvnB5xtmXaI1tobxBKJUVrinWsLnxbI4j2eUBMYrgW/p
01OGywVZCXiwvSBWJBQWLirkyGjjNl+K9w6L+UBEG4fNUsDVJchaI+XAvFVAwtkkq/isuLXs6EaC
/RHb8n9DBF1GRDCOJMIoUF5DSIrCO5d9GSsBfmX7r9ANHmjy1qNB3DnXLcoy2IWmLXQJRavQFsgS
KMpPE1yhJzdMV2B5n5KWIoBzrY5fn56F/8YlsgJV/1JAvNnXye/jE256MS64LjzXJZMRta9NPfOx
XQHRZfy2WUGtLDoqtewaODc7oiyd6ntB8x7mT4t+Lw+81gccVFK0eJfOodQANAgyBNPe4II6t3aE
ZlQsprIi/8jLK/Zx9wD9FkTZ/Kk2yN9fnqPY+F6HxyUWztoQOq9WpbA+ZOvjUa36zUwvG0IzrtPE
2pcO0HzwVj0GFHF+x5bgz3xBHSi7to1t/QNdNRhwVhBZGn6cIJaGWsotRM+bizzQYNdvLezeLi+Y
Bodf+DnbzQdFKi9BdSmlaYslNZLBOXJgFFOIDuh0USPuCfePlvNrnq0S7IbHY3UOZzCVRoSUFjFM
0L+GrtIGnFdzKQimloJ+taQbPIaLNiiL98WwzWNfy4yy42/wxrEQyrxmCp6P2fQfWgD7Vs887Wvj
sKY2Vwb4Dwz3BhVUnu0jEAH2d6ndLbENX4pM3sU6TaOjigmDs2TROE7T+x4YgEF31YoLoaW4D4M0
kluMMjNRmoeJAZdXLZ1BTHvp6/cfiYpK856+YoZqGUUqUZneaEmbg40WBhtDLthHp47gcISuyoNe
rYmTvMnpS6hSmRFA3ra9uS+YwE/yM0hFEzVsO9/WEMKm3M+hDifsqofSNayMmA/STWXnNkqC91Ft
hkz3yown/zNu4Pzwt54D/R+T5SW23RvlJUSdcWKjCHsgaUkpG9F4POsbBuQGU/hwbmxIIMNwelV1
QmCo+jnpp/9TAgdegedyVJlQ04ACbh1fqqkY7/m2vlZwnf51lZpFrLhjOOkyVwn0w7hh0Lkr3RO7
LicbIFo+7l4EfibwOrBY5tx26UVvR+4RwnPd3vqLEt1N90os4W/OKl6dEb1w4CEhO3R4LuCChGZs
nwtCR/FOC1etYFYk0Ew3A+q7G/uEAQnKEohGhqrvRPviEmMveq/qoVVs0ScrEbANQcn96v3kKC9F
mQMcmk3Y7IDNOrIFqNUfqdLUEHuKrP1EnL99uQvgo82XEzbzvVRrbtJvKozYx01b/o8+1jTHRwLy
y8/SbJ9hTTgcyHElW2F5U82itRJWSQ8HJMm0Gse+nJtaHii5+kK/LULX91uXMFfJD7LmEOl4LuT8
Qus6NEbw0QytwVG51yyui7X+jG5/31gSFS67mAMmNab6dG4P0pjDrZnTBK/U3O0A1PqmY1YaSHEH
V1sZvfpxI5x0b0OQFVlBKDJiYODa6rHD4mEoYeliSsL1K91y8+74koRAZEEzv+nKxPcULLdICQ2w
lsFaLbmqjXtJp17oPBtL0A+U3VqidaAxDUGf9U8ouqMghWvlvypWwiQtelkV9q6QumFEzR9eOCqC
V5HHBFNW6HZZHvwCeKzLp/9/lHvmhQJPyu/VouHziiBMDPTsa+dVVpIqHmxB74Wh1ClIVka2dn3X
xRf7qBagno/zDnOW4wnAQN/mGil+Uc13IX1ceUxRme4FsiBgADgmEz2FSOfr8TPnHuofDEyoaOuU
nZbZxpRIEX4yL2Nky4IQCUd6l9+S+YW3ZAB2Tgisw6akV2OYkw2I9z73JLudYCykyl3s5fiMTcwj
EBxgNFq9LC8jH2piR/5V6bBaelgqetr3PCFNKhz5MfPWAz4+6RKCqcKVmHlFwkbRytEAWoFKepWP
E4XOVveqW0Zv/phcGra9YIOV2P/9ANL9GjkuS/3XgwfYhqY+lLaEoKghjojnr8TcQEeAwWV4wimu
NglarguwaKB0rweGB7tnCCMdfKuf0m5cj8xUnGLNa/XDkPBxNsXTCRzhYbWg+wH12n9AwiXQroHO
nDwpa+HwJtBj2h/af12hq9lDJXUvipfXX/gfl3AeYZOmodxRdOSMS13kkl0DL441xirH6xsSa7Hg
31QdjV1x3rRrF+b41kpEsa5huXS4Nl3r6Kl5yQHFz+0GiozP3yr+MknoayR/u0oIHRkieaz2GJ9M
qUgyR8rPynL7i8wwgtGe6YtKuM7A1ApFFVbr7eTDg80iftiYCvz8hAKnvJtECrDbbz8hwozT9QEc
ivY2nQrNGUrau5y7RBQKuyl+iPdazhSBW5VfI0DEVgB9AIuZ6jlMWYs59kShGC/7SeF5cCHislBo
F8uJ4gEUHiF1/cS/POZw1cjIrWxx65tIpwO0zCZT8Uaob8/SnpZHsIO45KTLt4EMvV+LLDbBJ3b/
QMxEXE3tQcToS2oZ+DAWN/cFvwp0nbdy02dpi/kSeSkyMY9Cztyr5DgVVJekDShruDzSaUGGRo6/
HbjJRNOfTNXEw2JCK+D1SBEItfW0e/BnYLfrfml/Mvej8f1iv0+mgZdC218YcRQI0W46fO28Yn50
W62WZi90e6zRT/tXoyFkU5tr51FOeuz1sVk0prehhW82jpDWj7rtD0uwCMiCbu2yt9JH7zLTXD3l
2rtPjyCEZUE4BvgjO544kxJo7RJ4SeLVs4ScWxKsKjIuY/0VHx0s+EM0Sx+3vYKkK+DMHrdDJZD9
qk6beeD+O3GnKNIB8d+9Kr2DSkM3nP9MM7SeJigXaGsezVLxwcW+MlKjXEeGhNFoa9Jd0VZJ9V2i
nnYr0BWyASMJXMBYL5tIVl05d6XwIPhsvrQ1XhpwT+Uu9odLZs27SiEyrhYutXW61oobscheHNQ3
kPS7kCVXH67trfiWrkSwwCzKt/MqAxKX/I1YtX489gjzFOuBi1gkAezSMfpXSp9m9oOE4jIXhRDW
QB2gdU6IY6VQVIyyKVUULzGOjiHxG7Vqk8L8P7dDAvdQK8RgNDj2gTa8tmpldn0JzUMz1KyGiIQt
lS9tIsZCnjXkXB8HaOMrS4v22INIkPmefHrI40lq0ueWgr10j5s+hnf2rkWbxVW92+i8afXqYMGp
8Z954Fr8KpbI10auuDhADNEopqePTc2NuNlSM/ImLdd6XF2/25OU3I+ELOf/fm5lrI/EQOUJxONY
VqB/y5pzuE6rPfVD42l3bMkbKewWXnVA39AJ0BzKp+RjnR7KOjGLMg/tdA+a1ViEVKl32wjQxoWk
EIIYYmDCPZvlATo8ZwKaU2L9qw8775MNnMTgSNOoOKfqOUk0bU4xv3fbjLIrsZsGWDLxU4xph0sa
DzWMmaTLU4HuGnKja7c2nlS5DzbtMq4awhtQRppYhRtb8uCaY9LV/uA58Mwx9Ifqd+2eZ2qUwIga
XZzPCmKw8lHSTxCpmhge9JoegZcVqDtCdKAVapN9MKUZRW7LXOmPZ2KEf9x+CP7d2KTPTRdgjK8T
bt9PrerDrucLTqgEpzUFVA4uAhseuSoDEtYPOlWIUEjqhiwPNfZclPPaxArVA8V4f9RyD3FXCLJN
7LMO8KfJy1r3YDNZFWjBVIH7m90wFu9hPiqjr4hTlWtBfc3k/AxzS1R/lI3RFd9wlyILaHzW6DIR
yjO+hkzJdKFidpx6OFqlmm/qnUt434+nl7x85pw9UDpYSaIZ7AAS4hS62kBYbCCv1+JB1py3EzUt
C5U5gB/B9af/acE1T/CZ7CbXlzy2DhS8hqWHf2N3ijEXVRmPRCiLCg2ezZdi/2cSjyF5Vj0TfZvG
oUvBRL3l0fGbemalD0M8Fo4FlVwREt6Zm5B7lAHoLfmYlejlCLAkrcjQ4f59NzlNT6Uls3onsjmy
51FrjBmx1MXSnD+4RpKzGtIkktUAHwhhBP6w6csD8vtLnRWsbn1LLj5MlHciJTDcCLwt8jDfGG8R
FOJPzsp1dGrQveDJKSy4WWGdIkWyqmCcNNE9fkuEqyrve1NCAzLPlZO8m38UmuRPLyo4B9VBlnVm
fGQ8g/eSLZifu7DTHsJfoxrAHZhBndDIDAsEmNkuT2rMkf+dUGi9JImE/HD4aTUngySCMyxBBED9
5ib72JKkTzAJ2V8UacAGnjor9k3cFZWcOn/UfXmA7WHF+us89IXSo3iOErE3RkenV0DnET9bDgjk
rpE/Gso23O1EL9pyUY8tMlqw3BxB6yF683ZT8TIhs0EP0us8JWMNwV+p+wgpsZuucnQoj5giGEKH
c8fo683sz8SUiyMEaPzSE/c0eP5uJRnNXCrazcNr3hTuUjUUFUgHww0zhedQhODEhCSq71/KRaLx
kGJ4uD6DJhciug4FOP47UA67P2hCFsno+0k6whuigyCjxL7W+zF2xfYkWM4lIpA2XKTxyVsrVT0g
k8LBUxuDFyV8YKYmS4NvZ0YDaewRBzgstOKZugbPQ3E5iLMRBnOD5piWHRbJ/7kvZ4aV3tuOoGm4
NljXhicJC6K2oJSVVSKplcUgatwzsyrGnRlU6bBN4CvGC5bKcI07S0W7Y+RsZ2QxYL3dfbGacrCw
djsS3/1Ca9DHqgWIi101GXMAGUmmOdJEFrGxZ+NwluIGTAjeUnTIGVxlmfFbl63Y7x5052zsQFfp
pB+wPJlGXP5ynq/clZCrLD1Epmiym3yHANPDE0ypamtI9dHhdkRWb3RozZaeh6Jq11lzBGqopBm0
WjI59qsGReObPOqpmBQ48Kqcm6C/f2Zg5k0LpUlGqGMlBPr8+bC/cQtYLmr3MMbOqcZXR264saOj
7n1ds/ndTspXaRbVpjECnXPxMYFG7q71JAfJQpmePs9Q7iDGvI9kMQyTzGlWIoOvvZjL78HbmoS3
JqzXmQ1z+gtMVhsgBEv1cO7eP4GDyb9W4NYrnCxfXPSlYTCE9Znv2qDMgY4obmaEAc1BrI0sHQEt
cXsFBRKcKbhxFWSE89cZjt8gbpzxuN8k6WmmOF8KmNWYSZdSTViVVGZydBH0c17YJYxx4YVpCIDb
AD1wtK5fXjZYD5UNPQaIe7cjVV60zRvcVyFE7X0aAYYeFCFcC8/zAHfhZI7pVWSkFlGKhsO4n8BK
RR/ZtOWb9ovIEKQ8yPXLKHAkuprtT9KUR0l57/HykrjoaZSWf9lsJERr9OkLi97pwwZ89uZCz3m8
1sPudfRsCJ3FNXiMGkcFz/X90EubUhVFHmGfoEjEvZuJ6tHLqaP1wcGq1490LhgIK0wvInMMLdA6
lACIhsO+mTAe7pQiRxX0aZYdzurckAtBtcnRLMAJd1swagcurJ5N9PJ3t/fyXocMA5gbnceGL0IB
nqm8pF2f6gZgI62T82sTmp6x3HA01k+B6hJFoxmIBqTqApa7IMGf8DLx+v39Nnbo3WSorUkesSuZ
6ENvXrypAycVewoAh4eIizaA2s158H4CFnVSDae4GzrZHMpteRWO0oD5J82wvGb4HS/QDiki+i4L
79tUFk8fA1dYNw+oZoyicZVtQrpOQZIDKc6vbmHpQqDrjidbXW3XPqhBhfZGDWfFHUcK3hXZdF7C
RpsXVzzkHAEGA09dPa39c5UpbSDmcMWKZjmzyuOE91Rltv6G3Mu+w/lSmLw90nY4JzpyzQaER3p7
CZ+7+nJryXiVDoZWpbA+xRQxBVnzZekM3telS2XxOB6YRoHjLBOH8rzJ/BJNlhHFuzSj/yGmNwtG
KAZ7WYTellTwhQyDaFTi2jl9W9ekEC0MW93W+jVaGfbwRdNhUNLgr2YHi0uUMlJcukQYV+MwD3aO
6+EGX4VsSU5cNXR4Qcr7gz23KtTEFMtPD9nmmw+tzt6SgX8XZfxaBI98iOgIn3aMlHPi6Bi3DHvD
oo05oIRvx63p2xxE+rwD8yh2bqHHim4uAbhUi0O0DEt0WzSSBAl2pUoLgfwZFJj3+qpQvze+2NmO
0Y3bDD8VODdvG6yKefkFToj4SaI50kH/7kJrNFooyIq3cYbMzX593dbvAE0LNMI+VZ1kYES+4YT4
4RHihSmKsjXGVj7elKcnpbDQ9k/diI/CGhLZuGgArPpJKYlYFvxszYvHLQPIcMDruw4oEZ40hr0I
QO7M85RDyAlgyNj8F9xYIJOnpeFl0PotBB7BG27kmpSkE9zm6FoIGtw1ZlTO30wZGIcSjrHIyxvt
PFwG2FnT7o4RaYL91sTaGNPVmhuup4zWTBJW63j32DNWgnQrHEID2+m2HWD1wuO9UetA54e7I8ss
XdGx5xgJ1MRqyfkRtjrALjlzgsdaQX7F4h/V5blrw6bUUo1oFJoM5BhVLnhb/gGAmoM2GrAYZ9dD
PHALlHBowA6chZQYKQQ7++816YuzvYPoOzF0KcDutBiUrRyQzG/2IkjqonGoqAg6LDG/GRoWooEt
BRfti6IPHhydinJ/tGJIWW5OgADKf1zFWi6u5VTFzi9ZHp1clDuoijlOg2IfFDA/75DkMu+nGtzk
P2I6sXWKeMUg5t1gtOn0zZ+6Gn5ktJHfLYnxtjqZC8mxuuC7gPEhHx2s7tBavA8B5tezL1gjZqkY
T0AYU/fVcTLk+TcmbQhvPwTZ5txXp32Or1HTkIz6m7l61vH002g8Z/avJU2DmqW4QW4fO610LMST
/7VHdaJUaXFfL/gv1nMR9vpAhqfsWH2vFr4GOBJ2x6iAzn5LkjEe9ADKv3C8ugJQ4HMLHBiDfh8T
dsxemEEY9Dzr5AtPNa1eIKKE3uJeCJx2v6erlCy/4dLRqdCr6E94VqTbRYP3WEF+dCXcV6Mzszfx
rs80zPKvDpahWhTyc+ru3MJNdLf/HRzluUPHOq3IW6tlg6WhmmweQxRJYvqDKEYZ4gHCgytnlC5T
MexhqoxMGn7m4C0bXAdXWYkrgjXpWo7AyiWLaJ1qwGZNjAeAUyLJdF/JCo4Xdj0YMZacUZrjrjjE
NjLUgEpi0ui843qJ2O4SchOv4hEw5Y7GognQmrkm/oV/L+CU/b4NKYaJcT2ZTnbgWkZY5FndCSze
j6AnyP5nJq3JyFxzNtJMOE6xWgFkpC9oeWWSPlJS/ZgrAiRl+FkynMO/NqL3TNPuo7LjvQRsMZqO
FgETzP0MgCT0y3CdGGx26V9PD2eGuPy8saPyt7ynwlPINyThWX9artDxoDwTojBHZ7r8UlmuIhh3
SM8stPKo2KDbtwcSKhRf1WlAySQxVBsjRno4XkopQSwjtIX5Y15NinntDbsZoqySg0uqPINxI59s
zQT7XTL6Cwif7WGuP3iGwcHbHEPkEHnxaAB6QUy9ZFqiwhRi+oG7mV6qvpKudy2iX6zR1Om60kT8
97g9g4iUfitYf3L0Br+o23r28QK3fVm4K8WM9eanHiAcArGXvRMwyyTGQzlhm+CR18/6FDzVzs7c
puEHuorS1z5l82vkTDNqW90a+bTK2f5tMjgQJPF+xfXAQ+UZ9P8tBtYEmRLZe3j9740KlgO77G3R
T9jBmln3W43kfN383vBHgtfdOgZpu5go5eywShfQ4SYtpzCrHKoGeRRQ/Pv5enIQHc53uTYyOhfx
BtGZmQ9wGZkCXFxj2vCiDF1okgp5sGAVUb3NXzQy4f7zsYrxJr/2MwCwxVvFTOAqL5d+u+SEZBbj
VDhTC9nXZwF7kuf9cTARrH5qdzHJmlsZSzriViXh9zn21WNw4GqrEQwf6xJ/WSWiWA7U0DSSZpmz
rO7ta1M1VAc0257xesc11ep0nwD+z389X1ev1k6l0HgrDNj5GriXQ9oRDmYt2RSEeRcjgd72tUqH
5F6uKeizoAuZ/MaKjN5LN2nb2d4jVLaxKVybUq0EP9hLtoJyfYS4yzYEc95yN9EL1Z8S6wYYnkAy
vdAFvnCTDc4ZFlmnwK4H3fS+BmANBAluEwn9SeSgoQM9esfQYkrubeeKH2ibSzUAaqK7P0XNmuWp
zWks+IiqkaCY4XqEDAdW03S8mMPuqAvgsMIpmhrTcD0RXyiaa4WqdSTuwrrbWs5j/8jzhyrnOnxb
Km+ONGMeCsDZ+SpkhqdwT4vTb1uzbVOxzd6bOQQyBLtZVSUMDL3U1ujiI7DHKyAxc0aUF2/Oazx5
OBJemi7ZQVinNVD50l/PRGQiOu8b2U8953RzgrBYKMrSijD9ERttdmx7mYVv6v4afnKVYpAZ18m6
k2MCmzKmiZVT0d+2KJaZqT4gHsbWsVc5deiWF2k9j+adaTD62V57Zc9fzNZLx1jrEqBYT1C4GmH9
phC55HiDV7My1u4DH7cGBGn0t3wmu8IkWMpQ5V2UmbaMXP42ufBf7xlH4ghZlhO4tpePO55Zp+gz
RX9j1mQqxrwytbstFDPabSCZqfIvAJ0VGwDqgkbjyT9vXHj0PhSr68UyR4pwotROL33RJZTuZa6t
E23mTMa5tQt0yxhSV6Li5UdKg9gM4U54XAvKi5lgtJVsw7dfiPtMA9axJxdPr1IeLSHRQCKuZ6sU
HOmJmx1IEsaAUKlygsxz5pItkrcbRbtvWy9++e9qFe8pxPdnHwwghp2IB7n/vp6312T5OV0QXD0u
jVTWh+9rw40oLZMjdf9hEeKCmwkw0oMLf+713bObsy2vvIPVfoieYH0CxZ3/kZ/eTLX8kgHI6eWQ
DtLzV9Bh/JIRIhKgchRt9cuHrUhH+XnWdiAhMXrhPsJtrcTNw7div2Lhzm3VuTWnmO/czyjBQkkv
wjCytoBBvoX+1f45bP+o7PUBT60iUTcLUViG9RkW1k4FtJpNiNX5nQlV4J4Zmgl9FIWho1tOwBsI
kLnJ0UxTaG8zFl6hDkK93Grh8emgZO2l7KjmW+X9iBIFMagnSZsCI+ib34a16yIFpDCbK2/BWhZK
NUCmmSnAStf3i6WZTO2RFCbZOi1oFb7EbLm2HbZ3cbO4RjQf4TE5mEOrWGxsJKe38s53YkNUbP4h
n1Zr7438VjKh4Y++4Sc6O9/x1E4foq3ZDtwSMihPAUJMQ6/xg/WL0HB/1UCr7UnopJqiPx/VQepi
ZyyIvHKvDqAvIYyNC9Psff2Mpq6srM2VwNWAu56IisbO8Xx6FBxx9JNYUg23nQefHaz8QQ7Ab46e
0gq3mtq+ZFuzfllx8Qp8hoyia9MAvWEEF5ehGVs1n84LGmL+PptQNkLhXvdX9vWXGFPue1gWSPlX
RWswTHQaQd8xahKbcwCMn5zirkWjboLJ1Knw4r4Zm2ONoq+XgtdLGBty6OXJ8JG1imr79b+TOWK5
zqmK17DibHLGJphtODk9iJJ1W5LOm/tWY/l61gjjHLEJgp+hSJl3QZ5L8xou74dBCwrrNlfxrlmk
0DN8RPFemp1TFIDRphLiuTufMq0QA3JspzyIN0m9iDxbNnf/WBp/QmuiCG41DUaoDXG2dYVPTl5n
6FnQPSsFrpnpVllpm9whg/hxSdZcpyJMTjuB0nA7pM83Pv2mGL8OBZw7L7uGAs1kDbPoa+ARW+cb
HGLHLgH2VPgH8EvKuvvdYs3y/osYiLi+K9u37odoCJ1V61dGgqo/CPdtUZLzxvmdF4gBq+wJVhez
aqNE6SALELwrduC/mSKlC03neiWhwrTmwgX2PjW7aZGmDTkuumAntzQyx6ayxKwXs+atZUxzBp73
/0onVfjfpt44XhFih9SLAqQM2e+jdJu95sg9YI37c5tl8rtUOqCOWmFIKlnBZ4bF1hOmalKkCCr6
tI6/4+oN6okiwHaHdxJQH/Qa/dhPjMrA2RNwkTBPtT3C7wfi90F1peYGNXeKrz9kFMt5lwXSMYlC
VT64ysVo0px6JVjsNUPYPZk3wDSfsVZoMmdHbp3JNuMfffPqPKbPjRJiYGs9aNXaJHHzqQRIGUGa
/KI8rpdBO+iyHtRjAw7s0Z71X0Cm2HlantX/Cqh/aKseeK2Cz9NopP3M2P6KFhZPpuKXC/MeFwjs
BTOirv1A2svMBG0DK7ELJNw0UXvL8AI9OkHIU+PeVh7R3hugGSS4sWxMM6LNHBaryFL+yOy+aJU0
Az+MsPD2diQX3JwmaVfC5dK0eaNpco07zQvUueObxSGWQlDPyuq75KIyTgOkxV2KzEez7n0KqNLa
BPt4oeSb6q3itVqV1t9xce+FXFSANvWSC4+6askz+KD606jRMjI/59AFMoOq1wTOdZyzCMd/SEm0
Beg7rYqYQGVqQaRlnMXDv22gErp1DI0T3hSnSPnPQQef4ByOg5dmD15y0V8ETKkGqNS3hf9g11PH
nEW0iin+tCgl1Dh5XofMeDRjJcNIdMrd0qmNLyXwEAi6RpPUx3z7fTuJNbCtANLaPhu/oJR+a6Gx
AQBauu1Sj7x2DSMhHUuDAKeLEZimcJDFV8+CkSgN9m2Np9zgmCTQ5V6eokcnuqf/ZltE4J5wba6T
/3uT+f4TiWTwo2vfo6+tHvTRNqR6psM5k6Gus5xte7vklrDygghMDLeYp3ZuEkYVajEfLy6wlkFR
LMJxpHU26GuyhnScgHzcab/tjYbVc2bX1q6j322bShNFcTZP8+RlxAvH6J5gE7pcsV44ox9QTmq4
pXzMF+eHqRYmAtp0ogHqMDrSda+A+moiGl6zYp1VDpJUWzCP9dpU7F1JT1nTKe2skJOvb1yEpTny
SPZ5kG/2aaFek8h/yBldTZ1IcwW324qJEzFv+R34IzBYt3u0xPv6IBMi4e9stJ4DFRYflj9UKgQ7
Q/nQfgw0qSlUrOvH6IsdirkQtkxpt5EjWTS8x1BArSWm3puZ13H38/jJ0ub4bScJi5z26wzxMqq1
Wy7mjpKYu565ZjT39Cq7nLrj9VZvXlk7JRLDRgyIsyND8Jj8uUVha2fKOwojmoTA8p2wfSYX5g8R
2ha5Sbv263dBTJLDE+BKGsREtJ3sY6Q15zJbCmiZWYJsMhBo5HxZyhtOEtwJPq54Wv4BYx2c+ClH
YN3TwhGlOUfFCaIcVjd7R552010ZMdrhmaya+5rzjd+JDGyQBhyn6U365hQQl5P/jqgYfVB46Nx7
/IcrRPX7+wvIi60szOIu0Tbbe1PDwCj52SX2L765BpdrPb1W7zQ/XcgT36mGxtNNsgbcTlvcSfgJ
CxRtmrPaO98OVaowI8Bj4PEug8366bjwOuDovdoeDr9ql93IHL4wzhOAeWRPMSE6kI7gnqhk2U+c
k1rl77FBsTx0kTRIFaeFLCV7sMcAupPjF1eJNXrLHqa85f+FpYc4Mt97jPtiYjRDLkYHnmlSZJRv
r9cRcl0jDcQpWnEM+xBzUo+Uzpss6T7uA7qjuRXud/DwB0g6uNWEXfq8Aj9owhFravD+RLMUOSpV
tqb8xuvyj3xWNEGBd0EalDffoKQBB5FK3qXsPEdu3xaOiBD6oFdMKKdJVS8BHMXaSFwEMjtWVlzp
x/wV1SRp3l4z/kwL3dn6ddPQzA0bmszGHBY9vZ9hQdW0KL8Diq4VNQ/lZKdufwT1z0AETUAVcFsX
/7uuieYBHNAiY6i/aVRmVZ9QvOZxWt/WBzcpCKwgJ31QJZlSN/FO5/z39G25i0bqmluBTjEfITzH
I4nv3Vn0njejGRA1Zo4Q4dtxFXtUWYh3jD5Yak+5e7arpCAPBLRLb6Ss0uFcPB+PzNNumjRjiSPh
Fv2sWlRd7Rj13HaRsoEnCRyrlbfxSd3JaRz/JG/5JdzNnhsRky5gbJFb3tlZS9CVcnyJVC/YC4+e
v9nuvYulh2nIgQZL5u8CmQIrBFgnwGTf7aQq7qi/HyG4W5X3M7CI56xheMfXmT09PtO/tOsLLRrN
uvPhJ+Mya3MHHAqUGSSaFHmIBm1/QHXPzcg59XFwD/92Bo7nkXd2UF8KH/gUnIgax0cruWKPiVvb
4sH0xzS61TUKMOauuLsJOFepDUQXGUbBDtMSdQ9P3q7T157jHVzcAQItvILh+k+SZMeZlkehio2h
/xzvKjDK6g8QNyZaUNRzRhJ5c8tWaZLca+hOW9i+S+F3efIoCmhP+SVuCdQ9n6z4N9mfoxSgFxuf
XgKfXQ39QrKCiDfxLsew3jGF5uW1Aw8r3nnTb/pCP48CelbrTYUJFjlGXy0fO6iaLP0LYKBWUzzi
He9XJwSHrdw75RlZ9+7wQSRoguHbAxNDKnl59ukMNQxHqNtlEN4VwkRJN0IoLZjAfd8ZApPf5rOy
jO8SxSPD3Bz5dEbAoVyQa7amuGxYgCf+I24H4YGvC2jCOFIHWZw9zX+nz7W3mQZ2imPUw3AHWgLj
CmNHDKbQbrZqbDgn8R6qtzqgpYycblvJpv/M/Q1tiIZzjqKQxg5q7eBKPpfNACzWXH47aSOJ4jiW
6lGP5OovztchVrv26X15yMWX8xgo0A7c2F/fj1ufymzyV1YPTFLshyIFCbSSi7kcz1CItWKMzsFR
fx3VM4yFJM2aaOeMAXFRyYn9RZSsjWpr+eLpUN3bYWsLg0QSqnjeMD9Fuy7UFxqdQVhKuWzYLXwR
R/OVKoiz0pXxY27DbHOotbSyY2vmeQ1b2l7hfN87nm8CPL2PyCYhVHehTzrbUnmFSS1pM73Q69Ka
bkyN/4gx1kVvzlGW+Kok83t5zzrBk4mZqF4l+mWFm3HsrLVBJaFEBmj9RCF0JCOwJWbN6DpjKux3
IhhoDhmcSYTd0DmxPWfILRJIf/jPE7lpcG8bJ+e2Q58dpe/TPI394/Pli4WRRXhz+YqTIhwblwev
LQvNs0nNIdewwOcuXi4lBY0iP+k7gEZnpTCDvW6Ya2r0c2j+iUUQ7Jgo6ovCvPsAEp6jUfyWyhyW
zt0C9oCgWWDadkmzWrpjb2ZQflbh+l52tYwd/VTrdhfGGgDI1s06cKe8u54YbllcviA6pX9fmfPw
vCfnIq2ekezr9mKo8vv1KUlwUEigQBOI7YyYBiP8ia/MwrvOFE6FctLkg3gCnLy/d7zWg1c2KOMG
mBfoQZ5ZnRqA7L4qStFOqvy52ObohXs77QcKDencd3lENJcAcnIPo+oldRUOYcNm/+daqRm7lJmb
Q+mU3G8ILIzJkFrJM59hMg6wGQS+8iprfA+YpGveUBS08/2u2IHasWra4OWeASAMh8kEbFVK5G64
BIgach87t3vM7qBmt+ctai5aKOrsN6gI/KMr00hcCI+yuuqLXl7OvuTMAW4aL0bcbVYvucCWCwXp
rCrLAmvGZ+3cr0RPrR82X21utoKHX1JNOMh+XNEE3QT8UvbAc0Wrn/Dr0Iu4YDDmQEVx0nX5DAbC
sn7GX6dCHwGjTFRazJWzlIe+tpSMuTA2IN36CO35akMOIKBxgl1YxTj8Ft7XukeIyKZcybOmXMKs
Dd17ktwROLPzHliNL65EA/9CZ9+xSNqvL9duQysFtdLxJI3Rzd97hOBdZT3lV5mOzxRq8q7objQM
Xl8rG4CFW3dNNVOUlW7EFQ6dS0FcmTkbz7uMApWWWQ8mbHLAzxS51bs931DfXM69CIAKx3sXBvHn
oAmdxJNmWEB7uBBNus2hCzvw6UJ1tNMs8zOEuvUqlRWgFwKlKquSw2+t5IEWF3qZGeBIIKUW+FU9
T6s83NKMsOqtqFYzeUlAjqqHm1tEzwP6IeXmpBNqLJVNfSX3Z5yinIkpdWH8zVvuVJs4YCFo7bcz
eR0yMdzRHQDnQfqwFma/Uxl7KZIzxNAxLsKGw/y+a78zXBLigpBH1OCU8kN3b/tKLmfl+sbRbHkZ
pPYFYWgP6283f6fDd4dOwp65X7pVdjUQNdnPqj0ftyeORi7QPRvcjNbgYKlqIAoZRWWwS46QStkY
9SGx5nNBjptVYI+5f5lNMtjGBHoLyJFJ20uUie9KE+VhLWoCl8DwVot2V/Fa9tG4qGPfpZlUm+KD
0VpJV3rGkyUEDJJwz2J9UQ3qYrO/KlCnJCMZiIfzow/clqSVhIx/qEjUw5JZ1BO4o5ND9IDUvxmr
Z3p6vFaLkpa0+BR5MHtIMsuSvmYC/TwUjuRG4khTrbjDWrLNkNhQQohXESBxKksYbdcvnOJY4tpM
lOBbLfpbmZcdNXzjHKETjsK7g2y1bdMPpuml8GdUjno9tp0MMNBQGB1pubdOazRL3x9J6LdiXIJU
gLmuNHLt5uO2HoyDKdibr+1xJInEzNbVClX35RRu9M9n9v5wlsIj/0RXuNLLidIzAxQZ7nl62eWd
EgoQmKCqIqfarPnTDxQZbpkwJ5KZYTdDbHCCzGCtNDOG/X68chu8RAcpvqFa7uZgUXQs+5pRpRML
DHt49kl1XabMO2yqTvbH9+4m9tCcM0aURt+AaHUZfCPA6Rw7Fun5SVWWwL3jNNmSngry3eelpbeC
n/KOAKnIkgj/7Q7wdIAeHI/pl5CKTKuT/t6E/H0IpQ1En+0ckR7xnCgX/DvQTQx1pK3pvOuectAl
nlMfEQJMehxabMj2jfuB/0K2/u2OhXIIsd37qqkLyPOUhkRB8y2a4VPad9JYsgHPB6d0S8Ntz/CZ
vq/atYyjL6bz/c88Kq95HR64wXQ69KsGXdMMWT/Oi+yvkyCxodyxLue2cnLdin3hOQJUGkvsKKIL
L20SYxsL0Z5wnXz2VuSfSUBe6Gpt6M0J1pmwv5QkebTYcuJlxTf6OCEZmhZjPiBOgdLtdsVZVwh+
9jHVzEfoGsmgQ9nAgaQWg4Lh4YtlpksxL6OQM1unSsdF78/Q8Tf0AV2huzM60GASgBxwT8hcItT4
circW+vJctMBavS69ntW3DfKADse9rFlOMWnwVnyPsW8+RhwUlE6hqRmtOznNz3QtDW1t4Xvsdss
gzs9upXspav24BBYY6ZWNHFzIG2is/wVmdbMXy78YaNlyYLyszA6eDT/vvHywWZBsUhG2q/Krd8t
akG6ytl+YdTA12XmyMe+Q5quVXz6UNwqybtcez4dYkvUeBA7fo6tX2HesSd/xZtAeZ0iE6wvbIwm
xJZ0yAy4kb0hzskytTWCgiGuD9yyH8QFIl2ejt5omR+Ht9CMw/flGnWkKlCZSTY1MQhUUWcSuNl0
75SZCakU1V6jPT1eevVel26IcDJZbirWfqVQqKD/yU6bHO6C8hZWMADeiZnznLcW/pnVHB5g9qZ7
9/bM/YmKT0q2iWA8/1zfhm2u7NLWginYPflGZJlO4dUu31knGE52VSyJqgaqIh828FI4GBfxfIkL
HqZHvdEK5lJ3ixuiSubmKi0zdQmguJy1bEpjSzks8csMjG0GiQqjInzyJSwcOjAqVgLlPZdHxrPY
pTXf5OROuUowQ7qx7oRSE+um1jyt8jXDipJvqlUyQ6OeIvIP58mzPhujJQtJoIRuLd0RAKlP57Nr
CmLbWAdo8YZy9PPpe1ovtCb4KYY9YFuiFr1VhtgFznD3ZvrnmE1vS+TOiVHd2v5u9PAK6k/xCfTN
2ct8J3Uy9oAQio0iLHA7+Ph52JFhaFv1YZs/U18G/T9PiPQMGlmCDmix5ejeG9KL7Lqb4u6kN0OR
mCqZg/oGsGcnsdRwTeD2QORxqu02G2h5D+6EJsWPcX6vAnOUL9e/V0u+ABCje+Wo7PVPx0cQNbxo
gOkfyRO2qbKeze4TiQPW65oWXraeCq20JQV5ZnK57GUFXvDotEqfQHqB52/i4aSIZk74euomSGo8
CkUjrSNvuMAi0CJyzkVbHpN6HHduUvZfsYSl5xBAZH0ag0Xa4g196j49zL0RPsLAM6rxBlnyIUXW
toeSjCZhRdn49dkQlIfTOvGZJlR1ZoFBEDz99YA/HJysMnpPeEtkicxyJmyuOoGj6OfRLY4qkN1q
hkujWsVOYlmxZxMDaG16p9t+VqRpEbzqb4t6diGFfDWpsgq3+VjTUOZ1s4iVEURKgBRDJMavvoyU
5VgwXbbFizxfemfASbMg6eRTKrWKeRLSiahPD8mDw3jODtXbbpoWoyzJqzKC+/UlfT+DfdOzxfsz
elmrNlwSO7f9JdkC0rYs41SBBP1jh17ITkLONU7fFFqu2f/gNpLr92lg8zu6JJHgOyRTIZUwXA7n
JUc8rqzR2yFHBVNfR2d2WGHrVf8eRFaz6lN9kIdqjQVYsxvyLyNsKihDZUbcqj6po71rYN5yirlM
JUBWblZGn7k5f2802OfHKHwgR+ppG5yHL5ouZqFEWuSfbHuMpddZdi0D8G6yzk4V6+Z2kiaA3FCW
4s5nLvEvrXO6LAujY51BbGA5ZhfS3VwymRCn9sAPoBmjkuJMAzHO32rlYaPafQEb24n3nYdIAOl7
30tm8LGYF4qrju9NUU29gJQlFtDp/FE5i9MB7w6kWacz2A3dcB/xEUT1Hsx8TLAGJ6GC/DOL2Twn
lx8qvtNmFuUt/s0de0x+1IUVdSx0CBZTnd77XOKtmGQSEFEdLKrZTIan/0VcZEgXaSt+8JfCuDi/
5brwjs4VZqJsLUqrF1mLLLc0SX5OHi5y0jh7r30SrZpBgOL2jwnipf0Txm8o1hk2hOCrVaka92QL
QuG3TAQKcCcWNCmt0LGEq1wAlmoYN2c4Tf5ocxBX7EIJEQC7DzZDm7Rjjo8wmTHdbQXtarWipHL2
sQqeyjTXGGwjXrsFVYlCO03FoE+knuUOqQf0mcMMcNANfhqAbcHfIKrjprUOKlg5r3xWcGbjwHQH
GRTRV9EVtLc5vo0lzFsxqRbDPKB8r6wsJNiwJSslqCPqj9bDRT7CXdmuMUYxhGJXhu/a7WEVjoPU
ascOtUQzWmCkCdwGkO+r8G8GNWdcWuSykm05lyUYdXY8AxH2XIfYtadBp6dsD3hdylRMs1WifmdQ
wNQsg8LfgSHFbFlyBCOImov550Pvv+3+jvL11wLQXskLhDpNCkxHCd3mub1gbccQPrCnjMwhewCu
0Oek0yXQ7L+hNaL2Wc4wpUnR32ixIjp9v0U9TUxipaImezXFv4lErcUDKgNzhd/0DTFUmsACe8Va
xXqCZKrUWNzH4qiGAHP/6otb48yo3HJQ2Z01al2xHDHS0OWQkqLl6VRclrrI87nq9U5qYcwZIc3w
0kEhXZot+tXUoDFORO08k16iBi+jORa/VM31sJvvlP4CezeABjMw/rmTv68NdPxCAcgKk8lttYaR
/BPm6Pg3M8RXvqtKdi6IurI7bMJZXrt9WalQ4hoJJsAnX+uHa4oqXpVsMnN7PtAfGEtjCgVGDj33
f4zt+oe4QNRBPEAUWG8d+4AnfBrU+SSdbDtcqzMoMHp/UIK9y3+TrHCDUZyq3P/o0DEOFS2VPDMh
tuEI4gKQlPFeZ7/KxtYb8L1SE7eH0CfjwXyntBvDcEAHxFTJiVRrNf8kZLPVMPq56xJoy+W7qv+5
OgQA1EA2i3Vs2rvlxvJzLCK05hf1pNeBA3mbItbi84N1W86moBOx+dUdNNZKNugcr2fXne9WGgE0
DzDcNj9NX3LMNsg3gWgSZAmR8DfXvzCeHmavEXLHyEhRp8Npcgmg0l1tc8XF4o7auKhCJtrHABL/
LXGhFkgUG8/0QHu68+V3uFpBoI/tQMUzrHiSJRkPA3zINsQk0gEcCRhqciZ2VLshDPFuz7zjsg0z
uZ5opJ6PWEMAaQadiKqvoYv/CwBjatOFGiSBaiLh2fWIOJHqivvY8cK/PD2G/ojgiz2Ofo5G7UXc
rEe86rHbOQPVhmdXmGWs5aD9sqXUjPZwtC/5JfDjUUFaMNacH+9B/pceUE26Z53TT+3laA7Br5Ox
ilaMIUy4VZGoaL/dgIpwbgXXerGi2bD9IMHV21RHVMN4VVLezt0Owq1ulDoj4vlLO4kZMOT4oTJu
K9mej8aDtEy8nhp2jNQvNOUFkL/LHs4Q/LzH4I5gOyLod5rObnMAjHJJtoWu+wrAjjkTOyLBM+TP
wSG3tXwzaYt/KrJF1DVutXbv3uBlQ6OHS+c44G2SwMkgfvEOmiQjQxcpEalYuRxyB7NpEvmXZOh4
dv/N9iDHF4MavQ5YYltgvc2wat3KbxOMEA+DmF7TXCHlkob51FJJcAkduCJ0dC9oPSCDzReuENr/
7d+u7ZTDj0ki+b6MOMmM8Rwom+Vd8AzW/Eplzr90CCk8pdLrhGcDPvMIF5iJTVtJ68hbaSxlpdKZ
JPQjZc4e3SB5+UHFeUV9SAMelx0vx2RksXBC0Vgt7YGMi7TTZfbO2/MwS/N+SYu2JvyajV3Sk9IN
KtRz9mnPCObjenqIDKQjPQ1EGk6RBstfaOajEZyc0pmnY63G1/5E50FF0dL/KwU4ttwSeMkwRsDJ
u03XGhELlHkAT0b2jZdDpQ6UsasfNgsTBXoelDg0coXM7EynrUPEdnTUG9o/6decPHzyy3h1oamz
BnLGCNOBFibw1f9mkbKVpqcFV9JVxxE/rI1MAzM9E+Cdzhez7+EKRhXYGYghDSsiLKahRZD2vz3R
tJdgkm+2bAGl0l3W6PPTlsrjvJiGmGWtrutuH6whPys5syTq7lFDyiO6qhuayXWyQ0mDDXYdNaI9
eqszVDFdVe93J0HTkHErloVUR8ytTaLGFDi/WzoaOoyXjleeIlSiahbMRqitM60Bt5hO5t4NG7/f
Ii3wu0ANvaKVfsLpykbE2V6AN5tVe9TkJKFEdW6xkc/g9OZ5CSwXc7s3mDOUBpUz0YBnspD9glCg
2fP231N/sunZM16IN18DDUqKW1eiUNTmog4OQ/uMtPNHsaCPYTcgiyZmhQFqHPX/ImqeypgASBYX
QJ4Sa4kHMj6eYAYKztqQn3EOcDd4CgmeWPlado7IDzfXN0aUmfFQvIZQ7tQCnQO9V9ELzvZ4jSLO
Fjm7IpVDuD32xolj/8OQduB4SYRqp8Dywr5pBIUA8dMGNpaD7NIPaxqJmh0hqQYJV/XSkulTjXQu
AlAI3gfdd2t57BVL6h1WGBIhE+hwmS/+Y1LuH8B4+cFkjCO8LjS90TVpzu6joRihQZ1qYy43ldtG
O+eHyyVzXjIbhsUxepwp1QmRqs6WVCBU6yYj21EYDjPGGUpIlwaH0YszWzLx083w1zxUlLc4K5w1
AmGOpGKxgwhsh/CGZmQvSCSYKLcI3yxfFtxr8XvKuKrcaHzXrMpIjQZhawBz6jSpIuhUzgso11c9
/S+9LpbwjqQ0SrCzcMZ/gn3D94TFQdhY68Pv8QBzM3+P8O4ghcUGJfrdl68PK+4tkOgNVPcTJEjp
LPqozE4cy+TjsTmv4erEchleQPJWaGGE13Z4ZerZ16UsV4Rk5keFm46qDeqCOpRlquZBHGgcbbMP
npLvnq5dOziFN+BRerXtl/FQXM0lunhLjGl/rRSiftEcuXqAMU2Xgk10DtSexwj7mxxQx25+ZBeI
1RmyXK31rmaenw/0Cdu6/PFmAihYOxRYtkzqi1YzrhjKmXqYxKYYa1UxkRq0cKHHBVGyOKuZ/JDk
QjLaxUPorPWR95ZtEDDttvy+UfF3BYG4Kv+0glJhNiKeVZv3GoSY9KxvwRJKpBKRN8dfmlngyLpb
QkFK/83vICVmfqJd7b5xtpHtVaY2BMbRoqFhRDURUMqISG9CJlM4MhF2vsEvykDmbzcMjtUXhPcm
FVCmS5P/xcUg8n4wRSuxiPSRl+O6GbX8+WyRxZgeoCQrYyOsmZt/pMqgjZy5WbPpDvGZ172SCGW2
Y8BLXtnhe+f+ZK86SpfmAiEGWCO3ewPiWMBybudruZP/KXcoVQ5vdiY6iOXIhSrCL4ojgwO/tauY
I/LnQZtmifj8qOtgBtaFpG2gXqGSfZr7fw2Y1/BOOEjyle5lHKXVN0bPg5UoY6gtyXm61/1qt2s4
qcs04gfDexmauPJl7hDyfp5C8VFxQpp0UWdbsawc6zxQ0C2Qa4e8Z2epP8mEA0ZSnBQWIH3936lT
tsrpQZN2EDvclbguA1WnuhQz+CfpKwT15rjvvoTDAYFhc2WUvFxO1lsa0MBfiJzvqP6F+bs6uhuN
FCwt3ZZn90I/SR+ZpFoEoZxjl2SC7yJltkQ8C6OfXwht/lIPUU7rOs/I7uCiCE6PGp9Sc5eAdZBg
sM4EIVjODirvSHmPV+uxLk91WaiB73mfEJHH/l+H6wG+iTZ0Fjb9tRyzSovlfo6nAPbXxYOvns7b
817ypocnPOSltvaMCHYZ0FMGopYj4O/SBWyKxpeP56LBbYlRefRMnL5T/lM81rXeh3J1fjRFBIYF
M8SGs/Bzl9qQHHQ/n4uHZNWiUI0nHrIW0Ttw/Q30KXBdeGoD1secLT7ZgqBv48DRmSVTAy8TURvu
6Vcv9oOL7qy1YaiCDF3MKaD3Vq5OUnKFsZstw5H1qyE/lwwD3TTfZlOhHQj/18ml4Sdqo1XRYukO
RHn32XpmkcgsDqrjqVIW5eNtVc9AiEYHGTfbHF7+nEo6yJ+txnYpj05/nGOYMSsKgEbdyD1MKALH
dQis/rvVz1uZ1gc1hOoBHIHRpDVHGt21Gmgngs0qOZ3EWOVpElHP5BQ3QbyjLdjL7Yw1oHjvgZQV
Kx2uGbltKKisE9SCY0z2HIT7GB3bnVsef54UN6K58/GzE7B2R9oZTSguP0G/KVGEwli4XJD/VXaG
6n8bJx0PcZ9/BqPiOZLSZCI+oUlTDxbbNNfV9ZQ7s1vDYzcStrCP948lobHb3QaVN4iaYRsnUWkA
0Rlw0cLqxAWEG+WBhbPzXaBC9dH/x0shaRRUL7kKqy+0bvWn+nFFDkgO29iFAwBKNBuhjpXgAQ83
9L66ZDpvRNShMFtqLZjRJHc0otQX6y1wv260MFzEFGSremdp6c5Ngs90LEap1ZHVYjmtzkIxCsoZ
pUSwAHkiVGTCnyM5Spu9YaQUkzKt/wBd2SskWUwm1nYvNjNjV42yJZXWXshadOSGbRmP21IwfSH4
dKIRjRoEexfKVNhWTd9kDkf7UWfCbqa88/6SMYrV1PZ12LHaiTrz0qmHKjmeNZVpgYkZqylA9TCm
lgYs15uuhQG+p456RcrwlTYYL90064OV+jEBULmgYl9ed4mKl0zaKGDMjcco80doKux1U9Bhqn/k
CuWwdTJlEGXnp2GQxJDhXZWfPVsrNSOgSDkzK/rXrg5cG20nhcZM09VhL8PDB+/pe91cvBwBmvIr
cqgFllHC+eq2lgtPZEQyd6nnKs1LAo/3mVnOLpWMEPP8Uvm4V6M8SA+nSKmK/AcXeM9az8SwA9iL
iT1SunHr/wCO6V79EN33TuzIXMqkvuZ6B+bCb1FKJYn1EnNo4RTThStoc/SDV7IrbJGjJ5Co7UzM
Gink8PgOGbctm7yvmPfCYcn/Pjpyxdi8jLMCQcRPvfe0jwdTsGdsnEjsv4suJ311HvyQl6T261bS
9BqY+/ZLQThAfrtBZ72zboMEgG2PBg6zQeB/9zz7fJ5VF8Ztl6KNW0IyezLO2xZk6BOVTju7PYR2
mU7Bs5LaxI7B4gm6RYSCW/4TubIhob0jEd6JOaDxyOXgkL6sXg2/phKPpo/D95SI3SLMXx4YQX0O
8PSymllIpFDyTWsPuAhzrZ3fXVQpBFa5ifiBzPCUN4r07MrPsBelNehm9nkkWHydRe+UZX5JbZ6g
IYMSFaNOsQ/3LfW7zcnKdesrwaV2pzyqC9NOKBnJOSUTVmpqnIDfniRRiXNIJH8IFgWscamBJShQ
fok7U4Cia0djQ0r7n2dRFO1smblVxsogV5cVjGrAE7RIvJ/aLb5CF04jjQwLcuKX+iZnImXsUV7o
xef0xV1z3h2Eb/asbzSM7ZmFSriSrbGILMAQo00q6a8c2pyvgU55iY+qYA+roqZqp0Dg0r347ies
K1uGDgtpuIVT+9MCbkTm0uQ4+9KUKIMmOTXnm8XqKW/i87kHosQ5dtAlKUB5+eKbSN7x7NAQxj+n
OE81ql7NV7H3O05QE6Wu8PDZUYJv+erkeIhtw7+Qd0vXbD9w+FDHTSrZdKhMh4Q3PP89eeOdWgNF
rzeMq6hRoovpBKBHQbBV/rhzDotJIIQv8MsVx/zfXdBFajuYxckRNvdIx1suTM1K9u5pSFAOQYfY
gLQq6YkepNPMeS2HA3FfUeYT4OAIRbIEsyh1ycuN8eLXq/SHTbqLs7UTwiWajMqvKNPkdxF8UMhE
xbvsYN4IDsItnEmRYJF0sWFDqVXqDaOJ9NK+KO1qBGLYlr3aHEbUKV9H1UzytLAbpe7S2Ny4lq6w
8fg9YrVTbtsZZ2Qod8Im9/kCj1ft3YF5EB09JaO4OAxlGAM98XpuN/zVqSW2CcsIhdh7jExnAyfx
MGs57hocT7lsPrtgyvRSUvTJ1eUhb7brY738ezq3lUUK8senF2E37T1JXjyi3uul+3TbymQ2C8Jn
DSoJIz86yvLOyT81s8Xj5LtqkXvvUzsACJ0e/EvUT3Uroucsc921SOKVruBiEAMX0dvhsqwh7e2S
nNh5IiV4JFGdzKJgg7t2R4gfMuKXVfohDRCR1bvnXVdU6tLQIZ9HrO5X4S5gw1GEYdWEFqZk1k3U
GdcFfVZpeIuc7u2vjtYsYgBre4TuXeba4xuZt671+a7UMCwJdlO4A4VB+H7sgffRl8VMTIHuC+jr
r3uTd6H1vdj0WvYzfuI3C/bzt4Qo/fCee359g8GlQeczCMLs57Ut+zhkSbTVTZOU8A+3bb1ZZX9V
tCVf98T7nEQOLmBtNlLyrPKKbIfn+Go1WW4dmkIe8WQzrJhRHkLc7eMFrBnfj77fbwj7aLS3+WbR
wVKJ1YVbIoyZn0vsCvNtRFr5ez1vLhBTt9BAazP08zdR+BVGa1hJjH+pk78Qc1HHsxAoeht7pgcT
mEQ0m9xCZkoMNi1whD266iu3+0V+vjI77vU/vCrM2cn988hFXMkm5V8GTcN3jZj4y8XTZh/uy1HD
4nBrjy1zlYXVUcyINITx124IO2w75qlh7AnjPCb06DrNzvgGAGzfv0DD2o4b49dAUI8G6RUUXkPS
0fZi9u3yBedfDdU1/61Ezj8iNkDratgY7dlrubpUkYqgbyrGgsrUJFWIOJgoHkIg5pI9V+HMFXzx
k2EkSVacCfn5a0QnMWOdiCpa4tUP1iAOwtvK6GcVf1mYODOO1cA/2zamkKphr2XI4Q/pEoW0KXTW
3TnpANwFNvp8uPWap+4MP5b8Q4oTGikTbTCBcZvNFNfBhXXTiRfD1KWX+GyESVx0Y0m2bPnHnSJw
HxiHSxGMm9skFGG/YEQdQasudgQs/sXO12Z1q3hCDmnuobJNiMfgviuzRgh09Ug7d4QlzFEbku04
Q5iNRLp64QxCBkc03fQB0Ywo4iyR8c1OCksssakxXWtO9Ga5R0WiMd/0efEnF4odJrtvIR0RCnL5
sjEpNO9Tn9UJ4wWdKpH5/W6dY/LalcwzucLH0EMNsLuloEWA1fwEdp4a//CHEFeJIe+6lBzm4azX
6GmAokr4ZgKVCxg7upURzSwLUUjh+4qdjxv+/uXvRucnIauEVBNpUt8/yU3SiSOZCBeJdFJQp+9f
H5bDqZXthYmyLN8OqIBgERycpvacpNnJYmYSiWymU3qpszlDdcDoWjVb09qMI/+Y3BlaNxLcaZLp
x4UEcJK0tbE+e7eUf+NrThj4Omu35Kvkcpig3dWOamWBBvL8xUxBmkHBUZ1PnVjgKDNwXbUyyLes
a6K5b7sczX3WzjePvwWYqjH06fLtFs5fM7eph209QIcaogZ93G9AZJbqFGZrASDWbXL66GWsb9fd
zF6g491Gjk1WHo8k9dDIvurFGkHW5ohwP/zUfzTNFWjFG9t9zZ/l1CFHBJUlK3cIorUs2FEnBhk9
py9SJmmWvJ/KJp3hAbLPSDBHctCnZLv57YWxjsf1AcuPDUC4WM/dStVlOcoPn9zP4Q4wS3QDhvLR
5WLpOuYAKdK9G0Hg38mrrA9FFzdp8iN1oEHFC6+rlOZPuTnDYdCB7RBb2244VuQjpzc907Ba5ste
yYgJ96Hz4z2JPAFR0+MNkmpY0wCk4iT5F8n9j+AFhjUZeKaI0P7PvzUIeLGQm1q6LDDsdKxifOxV
GUplz8C+sEyCRa8bLm+CSem/FbFaSN4FBPUVRE0mn2pLTS8f23SaOdCjiAoBNDvWK8x9FtB9SNnE
5vCTg6jHk9Nb1V7DIPWTY7PGNMjBnp/6i0WWwwKKd5MCVjXfrASC31hWgC5un1QLMAX1F06nxn6u
lDug5tXSPJZc4UnRYWzPMxrxUrvVaK4KzJRAMrg+wq/r8dAlf2pcEpCPONiGBSwLNnQdsDN/SGw0
SPlEYYKYPyRAwa+Ig6SRLOUvJcIg6PNK83ShYE1svv0MfrEeX6H1kXUYgE4TGxfyUNdWyVa2lihG
x+OQpi7XMPsJhSbrvO8QFqSHyF5E6Lzo++IF5tWS+/SW0rIG9/e+OaJWcjnfU2CnLHkmd1Cn5VEZ
SE4KcNzwgY4dUnpYpwdxIdvFA+oGAPloy9xcU4RXo/vseNNVllvFVfGyKqB9xuRqjI2NTPf3pqpZ
su9LRGM51Qi+8V26zVxTvRZw57wq5FNwG0dUnwNrLc8uS5R32ZMUjGYac3JC2PYM6keG5Iono5it
qkdagQ5TFK0EN9SNMH5f3Prw7ZoSGqy++apH1YCfrtuEgIZuewFohsaJZ4J0nubbtvsNlus0JO0Z
0hBPnI4B/jSgXPfvQ5i50YjyS7Pqs2QuNs5VjmqFG7aQNWC/AL+suYcHBjYkrEFKUVa8i/Q8cKFb
epvvlXuqZsqqNoPMZW7s53WZ5AurxafShf4DYE0PRy2IZm+rVWU0bx+nVLMfGYKAMVbsxKLn+mQK
/eDB/IAGAc5b/o5o0QYxh3VODLuIPtq3pOJjfVZn9SH7e9378J/XaoJtmtyzYxcXBRBYWpD/NqEP
6ZXqOwIT721BPsf+DYjRDU3M5uJ2mzLi7o/SkaUcMdc0AidAPo4trxkis/h3wPzYLbx12GLI0/TL
pGhut70k9YJS+45KQL8bJzZKJi7Es3Y5AI4FbUgWyoArt+qeFnWZFbHQ7I+EksL0CUxmFoL96srA
0etDDO0dIw7SusZAQCi5oL+fPg1W44yzEMpEc2KScXmp9XxNLeP0OhEbAsMzfPb4YX5B+ynCZtS6
hDUyaIkB+hHJPjvl8cnUkpTnpsIGEabGNXSlyxxnBJRUkBtRKN0yfOIH5vBMFAla8lbV3Pb+Tj6O
eyWb8sgou42ZyJ2pMZbBIi++8nQNqHFfLdDA7xC82vv9uQva64fuiKXY/BY/BYEIhHjfPw50hQH4
tPNnfe0CMqR5o1fWjR8+AezW5+jiiq2kF7OAdcus8ETqLb2Bv4yQN6bXGEkbJG0IbMRMhxxyFLyb
VsoNDtv2YDgAH6u5i3tPoULnbuw80VBlDPjT8/Z080tEPUoYtzDvjIlzveyePHVJq9kZJRdi5dP1
KfIVXfjO6jz9V9t/S8A4rxOv71tGJ3KKjH0Bqz838w9QBAznT08mvJJsXlbIsQfrjTaUFirTo6Q0
eEGlQxzF5CazMttNSCqMHRnsVkpkn762MP8pJqpiAPzaIdIJTI89iG6KJHjrLPNm2AEz8CZiijPX
/m3WVhbNfHIJLmLr4vWaCGtvCxx1oZvpgxZN2Rk/tbcXtoLRMH2LbbU9fOrkxKwR/qC8IQzLC20J
PEWgqTb32oGPft0qcVnyyj5fwKGu3S2gO3HqKUCs41TtS1OSQ1mypFymUbYu1nhpE7H4pU7CXvD6
uRLiegoerbVNsu9QqEoxudRdF5bffzMazCEpgrvpHT74api8Kp9ry+lH8rwO7N1VFFruyPm7T65y
HTuiZIYi1Zu6bKpEYZx1ckkfa76nW/geC1PF4VsdRxuiXjiQwhOW1ocDMtJy58ztxvIP4ypfNIRO
AsDo+1rmv1FziIvN/4vceKfsqLqySsBxsNV7+TLGDZywgYeVR8/rxGgH3xU6VtikBvAaR2JFL7/U
ijDmElTi7qhsxD2u/WNAeRTr6SS1ha9ShLy0jv/7unr77PokhKg6DZIUWAX3o1vKm+0WnnZTC7g0
xf1UATbhY8cVqtwP7kV5CJvoG5BV11sYTrKerhx87UKwpJeXew9JjCCQyAeI51z6/gP6K78deksm
E9URvO1HWhgyX/MFqPHeP9h9+Q0l0PnGJUOSOkrutskuaT3qp1b3zr+h9Fou9FUE9Sgw27c3fHdy
AwE/06VYqjh8W1DnWDLf2/D1fye6bPvXktHk+h+m1yOruCM5AE2U+2WfD2MvdwwA2ZpswsgS+T7x
rBXGYwi3MOMmnW6JZj+pBKt0TklROLRQSAiu1aawYGOzgoh+mBkVWNe/Cyth14oOMkYXIJGieYKY
PqupC4rceRRkc6d4CM9IqCpNfQhHvdjlJv+MhTbxpPyEqiqWVCOhssFlGub3D2afmYomnSuS4ek/
Kj26bAd47ejIXF40Y2frRby0CvcRgn9f9xCpErGTdRu/a17Oiyxc2cXzr4wXSh42KzR4KaZfxSmP
tsiS3igpbsCY8zT9B7JyzVE5r7Wb1irLJeEmg5+Ix2+hGIo/3G2wkcyk5gAoS4yV2XaCpNQnI8PS
SAQrQd/QkZIsobfdvLvtmctDVQi1DkLmtvTCVFUjaorf9EasAt7TDGZgz0mUerTRtqtiIwspHIS8
6o2R4yk0wizi9DwoxOWtz4Zx4DhxKTvOYlb5V1A8d8w/Zc8ZxDAjA9NUDYq2iZNodx+fNJ+3HHzp
3dj1wtvA+GsZ0uEly8s10405qIkrPwCHIDxN5ppnW5yyzSm6pi/taEG5KQ7WsFkIV/f/+92FX1da
MzTvN47cGqyJUmnMGPcCO3JrbAThg3HgWviH+YYRC4O4NStmz2sujRr2U0tNA6kslkR+rUkwSnh4
g4RVqklyki7bZMzcXy/Il3mO8kGeKCDxhZvuUeCDb+FK3VBsg3g3LFpX2GaC3Xxgx5zAxgr3HzUB
ZUMRAV13Ynr4sKkp65wJIH7aRHNO3Svp4m/FHr/KyPwor036d5/rPOa0otTuLLdpz4Hew0Ck06ye
ShIehWNHvcwwOoGtTJ1jBPfx0jFccx7jv++g+vseX/wA/bJoORJd8JdyCrSgCV+Z9Yg0Ww5oeyaa
b4EV8L1bu+ELwKygSAp1d9U8e3s1Qp0J6H6/KGEgTsYBhwOo+8MLOImiuKX5RhCeKTLGrHkktj1M
JgafbMs/Llpomtoch9+imwNgzbVI1miPUD4zY5sqBenm/aioLDh2cgu9Kh2BNRyOrNaia0kWmEGq
e8IEH2qqWUX4qnfx6xCWhn+nPB6mBL9LJBs1YDunUoHlHRr9jy/Wn+Helvpr64bkF7TC/rd0VTWg
dY444d1M8fe4U/V45u7PUvbibjG7pH1bYfrdLsGV3noaEY5RsqIp3nUOQUqszD97LUE90YBjOLaM
i6+8Nw8fUdN3fqnGn9tJL9+Qbyp9/a5xYeEV6XGzIpiuxZLJIT2U8c98ydCRG20hduIU/9s8MEmz
g89OHm7sTGvUP0Y5rF12qMg3vTfAiF+ehihVYb+t2GyQU0YRmYUq+dM0Usl52d+rQt5pVDe+HfyW
p3RyH1dLrpMpMJlt9NT+cijQ6rWiwZRvmWwOvdCE8itUjKYbV44nZxGhIRa9BEUNklxUNBPKxLch
hBPzyr3rGemhBpTpHvBBLc7tTzzvb8PG81lothEHv1+r5ryu+vuoFPlt5wCBYeUMLBsBP1zcTqp6
hSlozFNUYWwPaZjImrXR4H2gqAc2ZV2sn+KxTDFiTBD0tXt9R87v2YCYaujQtYFIE6LGTz9RN7vw
ZBw1xHvdURKljxw5IkIeYDnZxQYiozsRKmjmIyRGtKzx6FeAHP028AQkOMWP9CzoucwBcMVYSAAd
xYK4Rh7YQwbcVDuoYlfVNvAErH0BtWGPtwMbMUU6t9W1tGKSRYTblq4dQg4H92RyBY14quzsrsvf
Svh7V7hDI3uy5pS6aJvabXvwSOg/8TYmonNKAj6Z/VpB/OZn0hP94B1riKKJQGqfgfYsTb9E8Lk6
ITzfKyWO9XXXNUi6iS/ru763r2ClH9GRLlABpQ1AHULiMFVVBxLVn8zyH1JLLLecoSNUKXsAa9bu
aSDm+e2C73/2fX4b3T8zxuSmoNJx20wlB3lC3RmrOC2yqQU9lIHTjZQTqAgT2Zp4kxk2epZ5/SLS
EmYSCIUfs/7zU8nz4XuzSp5w6f/+m5nNhwl/6h1W1/jLmOxhb9iOIXd9yHCyAfHMRsA45It1yOY+
6/9qzNtYsSwu2jIG5IUoRtRS9EyMGNkaHQbFpSbR2lN37iJn4NseBZcvtY9hT46VlD1CfEB4jMyn
XoijLK/fUWXmiXOpWiqJbEsVmV/2UqlB0eXrR9HRGTltWTX1CKbHvW1mLE/N8PaUERGWAyzhnEPu
0UbKeJL0R2pdzOI6jNhaOQYW8/yQ4SWyLDvPUf/1fe4Yga+6pKtpxYLj7ax33gQjWVKyRTebt7bC
XsiBDVO2o/DjeorXlmHb/bjzIfNK19s8XEvBANYFzKKLJOGZGCpeBmb9FcqQO03Avv72GkCHyiwT
F80ln8Ph4rvk5Ycmkw4RaR1AIdg37gMHGPAcm/yJrBErOH8xModHgAj9LH15OxDZYJ69zgF5lOml
vVfFYVC0tHl6TLZEXjrRBoyBeH5DxDKZcltThvzDYgGA5iuOdL7GaIl/2yFiF73+gizW4SgKKYhv
Aqme8c1B09EQbSrlNCIDda/B2OM+bWDjfpzlsDKdzz3Qg8SIQG/5bYYHfnM60oe78Z/uoBkBWuHV
ZbeQ7wNDLfzQYMwyYX+exgsw49ouoegdy4KcFpCLf9aw05tluRyXpVk3uVlW4uzgAyodVFlbFRK5
sjEmN+iQ7VEDP0b4jc0F69EtcIHAvfywSXDtGz0iYJ+4TFjnYeiXTP9wfmskRxOt8L2Wn6fTuVuI
jRDPAJtDXMf18T6kUJNAx7gt78i6D8odVEf8tipASlz33eyXg9GlUxdG8neHA03PSEiEVVV+VEfP
zO2wN9KeprwMoF4CXza5iWDZu/BLXKXpg3bz2cDjdMcnP0cyvs7NCdlyKFaaSsY5u/tKotWO+Uzv
/U//FqcJWoMhiJ841ELDkzmGNNZ7ZS4iFLkWbTt0sqtecvJ4axhoY19G9HIZDroe94C7pK0wViHC
X/FgixpEHyw43kwvqQKN+VLudR/otx3LMkBtG2S5M1KvJXU5jEJbsGwVQ4u2P26YpPCRCvEs3ds1
iuWeKqCogxJAit3lxKS0qXdOVntsGi7sw//CUJf8ywOCyGgY05tFx0PClbzeQ9FyE8OheF9iET9U
G8GccFNK6SNPzDpUWjkpAPbpRr0uCWgRrVD5XwxgG5w3azV8kjqPjCLc4e1UyLmjqs7r73ru8jZ1
GM5ohPv4Fu+CYPOErYqalBBmS6K5Ui7YMfVexo9ZiRl+tJLH9scbmnkJWt/LLsQtfACJWsyT3Lc3
axM3cixdvKGJC+COg6WHShFJ46YWtiBeTKFPbYgcFT4dQA6bd4VK+4hNl7ZVXchjiKVukMqGe0SO
dMJdHtqWnxVRZEuS5GGdQmA1vP42g9fXA8PU71WirA3iwuFaxABpCnR8cS+KEUeNCBLpvxXiFip1
VXYgXEBm9ZX732ABe/eiqYFnN24ejGUlP/ZI8x1DjS2B/BJe3kMvpskE8wB+6Xl1ZokbqqEGcXzj
iSsHYwyscrJK3A13Vh8s94Kle6U1wZ9Wqz3yCqfHXE9knpDgXheaEhWwD5A+xtwfQuLTSfFQg/P6
bZ5tEzbW+n+wJM2vWPK9GsvMoaf/A5qNykK7k/BooVB/zBGrINKaR46vKimAvW223+iJyPGUJsfh
cbuqjRiB3Pv7jbKZpcVoIdSnD0tGwpLc6dp4BH1NtZ04yk5RmdVSnoWpZQ9cdujm0Whgj0ITIloW
wV1h+hb+vHdRDD3P6FvAGBFlVudKeQs64uwaSNNI50R/7xQxwcQISzLFEqhMYX84Ln5KRFByBfxj
JJPD5l6rL3B44TvZgwSytFW/agZOgCemJwQrxWgjFEgnXsIUIntuWf2Iam3AY1G5Q9fsm6uYzNFO
7+AFDlKO2pcvgyMIXejmBdIlSC2eJmyku94NV2eSn61IovSOmmfnUzndyAJLLzSHhWrObU+8Tdt3
fvuqpeIRVKl38CKxomCqd6erZ9pSKfx+j822dhD8RkW2ZkogUVZkokQPJtV39NnNqGuMujX6M3M0
LY65Wiu3iTq72mD2ybx+gPvL6OcORIMCUloD8zjzzP3hbFTY17GHRgT1JQx80z9l/5d+dzoeFuSa
kz/Jsm3uraUYy2KJ0n25fuacpvszRHBnN5g0pu/tLn+8fHRRAHt1fIZ+f47FG/ldgyGtbCis5Ay/
GllUSOcgLFvdY+UN54RETF6zZV6syI0MYWe992QjGkj/P24RGPdr5nKXvsmA4Su6LJFVomsX+BiD
dRVAMeg2KuP5Fo6JyhUa92jV112tgMdbz+CB0xjZDFNutWd7F1x5Lq9sx4RyLAZhqLM0+xqzkw1Y
eEBYZXnJtfJwHhdAuhapea3kvXsKdAyAXW1omR4sa1j53hX/UoOcAkdx12E58H8Q/SYAB2j+Zk2y
h6+fW+SZ7chyum5r1IRD08y1Or4xLY/IT90QRvmEu1INyMEHe4GsH/5TGqEy/L/LmhNHRgMqLBgp
vq93AfgeauvFNDa6ylqAvpAMcZ6EncrBR6v/NjUYQ2SyQvRIBvxOXxh8o5HqvCWidOLS9Qaw8W48
fuDtl+nogI3VMw/qvUC7mcpg422pPZT1COuRWraukXt4kFdLUDAVa/Kmf8Au6IopAV3azIQXH2Zk
tgYx/9g6wzhYlevZROk2tmOGIGz9FCTMs1e8hI/qGM6pbk4SwjFHcxaahtwSxvokdQF01sj1U33d
optrWukBPEB21P1EVOxoO9x7nOHxuS6rUauf2XLQmCViTqmQOIrxlenslzK7rqplP8vT9+cVu1Cg
Mk5XUffFoRDtlMK6D+4ewenQNP41oAQGgzBV3tGjDTk17rCoxbRhw3qG1xt/7Yx6xxPr8Ri5jXoE
/9dY0s+h7rtZArGC82U7yfvDkhkQJMkG59KaYi2aXNCKlFUk81EMBoNpV8IjDUYX3fr+J42CdMbV
Y4u74xHCMS7FQPSaTqr1b7dNLUBMEr0dswfCTCsk8a6DB6WDXQAHBUGhUObmhkxB/KhlEaNtDZQC
TGDYu+oOclE0vuEjVYHUJgDYFI1cV119aQRS5nzhKDgIbezZUbr5ja6CxG42dp32LrcfM3q0ZGTZ
SxbnzJ3cEUP7s2G+TfyfLPVh8/t5BFODMcILlULBdkkWBnwsq4p7YPPaHaT2v3st8+7Rpfqr9QfT
6y5FRJyDukQmXUqNA/lZLJj2STkQ2gEBZqFznUPogTvkEJO15peswBrYLNGYPGaS/F8eg49RBASR
92s4arGGEO3bKyuHdCSXgUpsQGnMP1EbR5XE1CTO+uM+bNtSk+Cy5X7peEP820pkbOrZo1BGw+WY
LBugVvO6zX0B9ZHcpeePzr647lQ8+yhpWk/fKgmqYO5UnXYD/QjFExEUb3TpibsCshuWFIgPy3hP
Nf4w4cINbAZ7kKbf87doD2hsYg/c6qOkuXGJx/SucjKyVI/Y2axwVB1yzQSKH8QhKGCf2/MXORD0
i9TZmZfQ3KLPSS/n2seW16111i8YUkhlEo9Hi+6Kv5ahqbVQRJObFZGVB/C2Zq+SjDZoZCme0uHt
W1qFJUc/d4LOdJmcO1e5AMQzLcj1ze9TMnn6MXPVOsvK4eQ1Lt+H2bavsIiXXKBAZRumdjBjcD9Q
enig6PgjS9JZ7/DvpIkd0EeboLh4Z3Qd9zcwABIIjymjoI57S+t3pMNreI6pdwuvvH0JWjP6CFX6
xUjQqSCxVIKte5QXNIhzlQE8XjI93kLvIvOp9obZ03OqCGYVz5VCy/LjXRROLoAp53Gjj10K2Cwh
l1QfnydAdfAcNDtuOPDR66DUKb5R54kXluUwkM9lTy5Ev3jC1/5A+gZAk59mpwvQcWXbkSxtTudS
pO7/56iNQtXXuaUcu2n2PEITevfl/6+BxqTULV1VE/EA3n4FhRO/tAXwk9BkB27D0M/PlEkHjkfh
7hP5mq2khkKRDBRTC92vMUnQdYhgLcpQ/ChmqkBU59mhJb52EcJNnc1TFoaLFXN/X7TxysdVaf3E
PwMRmBFZ1uolj10YBCz2emLKF2su40J/gyOaJ9gR7gsDqi33opEZny2dsdXT3coekMb6Hr5EL77v
UI4TvLBlkpOrNMrcb004nIQcN/Y8VQNaJ68cWGovdq9qJgnlvbj+v+goIaCsJuNHMzmWrZ/Fx3/3
2aK4KfSp+eDCXiP6OToJwlIOy61TkkJsQaX6AnEaUUU1SSyC3CUdkVxPurDxxNaHEjJjcxT73x4R
3+XOU7uvcLzJr0waxUqdk/Ha3/D90I3xHzrVw/iG8sbnsGXWo9Kk/hV4VNakZKFDexk2INnDWL3A
qs8GIRR2wulBV0MPq9hEGYpJ58LBXZoEZ9Ep5/cQw2xDuMWbjZdsz6YuYDBrhra41O9zvS3sQERF
zl/FcJUlZ3myXpi+ZNC1S0mVXop7e18zjLnTshzMLfKPQlcz2HMp1MOt/B9G+cnbFUfXhZthYE9J
D0al1waGShkYDnRQ1xtTL9a3KgRJ2eYil5UADgurHexhmaEj0VjzgWg7x61FrJQuJqweAJaZP+QW
6eGuj0WM/rkqB+gx37moS5YKRSTspZQpqPtRY8OfNecBXEQRpd0KF6/a+Ua1vtWBLmNDj9ltKB/b
ktGL4xzzFkvRNZ2vJ8/m5zUnN+W9d90iMK+7VvN2icX06/v/Cu8JOIGD7ZyJwM8CpwL+/p6BOlUF
Kbjrc5aEs9xJAfdfPM4ZgiPkjQ52ECOzkmjl7fZhqP/qxUNjO3nMD4frVXwn0CiIFjrAH6o2b2u5
k+273ZuZGQ31s5i0VIHrijKPxfjZG3rRR/hgnyke7KCq66Qk3bZ5sJQHF/3RYyJSgGeiPQt+j7nB
uKal9wUdS4RK/CFNyEhdEyr4/A11FU2dFEN3RZLztCNg94niHMtSGBEo4uiTuKoCy0kb1f/93/Ct
wcU0h+kcNPlGN0RKQZQm31v3Qai4iOc3DpveAgHX/mz4Pz8eL621P3dJo7Z7IV8HvbFI3C5p4wwa
0Vi83L0HIFo/BnA9ZD1d1OdBtSgONKnkmp9CJ+JXdKkBf984AjzP5VQUXdBcQvVHtjEN/44DVU0O
SAAewps8YtewK3bYzWoiiL88Thh8+CfavH+NEIq9jFwrSDoKY1aG4bnWRnCjSQekzwuG5O+Rqi1S
Y2gh2cLJ+I+UezEUzeDJAZJWfioN7hDks25tUMdprajuW3npmYKs3D5dMs71WtP6h4pTQlxIVaKT
3jufz6tI9TOTb1P53iFggyEKIgH4HhwddSHMKikrPsZgVqUwFaK/WsnRax7QtT9fF2PvncC3JIT+
sjzIrKKB3tPVGvgeHnusVEpIvW4c60Le26V48qzPjyINMFb+oWyMO8iBt9OQ/UXbBYC5dvX6Qthb
mOi4hX8zggYjp5Z155mybgt9hoklR9fDYDIPENCNRe8mbcKnlIynMWp/Wk5DVLgDvrfPs1+Hb60i
zfyzuzQmv7qa4DQBfIwHV4M4mGzX/9Ewh4EZyHu4vOoypszdaPPjRoBU6CZREuF2eQctxz2K/2ac
/LNNQDt27hbL01HT/DLsyi1DAlmzQYZhP/650jvJA06WCDnA0ICY4l/pHD9raN+icQJOO4iuyWfW
tZLwRAlMSH9iI5APszWRMHyTRnvMVU8CqQo7HjkBw0qb8i2KsqgM3hLo1cuWDGgY622kqTa5BA5p
llx+zTsTxxSR8KnzwI+6HV0qFQNjderd3VAOMj6adc7NU5lFjFKImLLIZbM4cd7oameSkPD7KtMC
iPNymLzuQ6SHfdeZQ2PvqFUt35A5EZagUG00p6jmkRUOyVIAJrFL+0MtHHMCAUyZT/6i7Xsua1ya
KvlezOCdqFms5+eOY9gwee1iA8KeaHEA4q5Moy/dv7PQZa3emoMV3RPzhh2a+6SwEpMuAoPkH5ZO
X3yIGVSxMUWVCEx7N9Eexr1T96hrnEnwlPIU8uxOVqhPpXWlLMb0fLUc5uUSxC8HthYvd+BqO37X
wC4K+HybiqfPwIzJ8oJ6zFkwXFEBYhX8haaSEtTybeBbjAV2bA8MQdTmDosp5cc6S6FlqWpfBa54
eq2yTGggW5a9vRaOEpp9reHlS2Zn/BJ6hkKvna4S5ACNl6KO4kf1hHeioFRl2P6DSj45E3kl5H7T
C1ClrkGX4FwybhbNmanw7E1gFxqJHnCk4AN1N+VUWkymH2IJiFCNP5z2wDUl64qCmZGiZ/am406/
8beT7R7njedilIKy2O9e40rO0OaeVbT6P+nxSHVaDzwOJ1EpUapRuc7Jedx1I9t5pr8/GkVVH8xC
ni6CyMGyPeKLYnerokI/yDZd/AN/xCy9j2a4B905yq3M8/24krqQSSl+iax84kgum1pXH0dVDwq0
CI4R2/oY7JHv+OyBGpLV4cvA5rJpOkXf1pFfOFIF9AO6Bx5hiiF87IJZGevBgcLdjv7zpcuTWhMA
0ZxEj6abLMMTHwxkDc4l64RSVPaJewTeb+TJeP6qycgwOUxMMZdFzkuHcBEuSvYF7yORuxGdWiw/
qLpKoycAjVNbsLnRoEBvtvoUIoxmB5NALvu7KedQ9qm1gMfK6OeAXeafriLCOmb0nIOL3dOpmhE4
bMJDMyd5SCTu+CuSukwCvowfXrAPVgcBWQ31OUJMeEyTWPK6znMR8FAHak3BAQlDSI1pnfojHNiU
wQ38EiSyaMQfV4yyyvkOi2geCrTaottpLvo5olmxKOB6CymC4pOvSt0/XRO9rI/W/BlF+4o6wnrq
PZQTZ4yMHGDqIaeBw8moYCBOqsCBVN6xZ5bivf9Rk4UpqsWvC85Lwu1+S1AQ6Xxv8E/cli4v78Zk
16FaAUk9M7ISRoSjTEFPSQvc+LSQVBulZyAzUL59Q+8GflaUzMBK45VhjMSK8zGMA1yisnI5XnU6
Ts4shiDuBDZR5wR0PTOf0jlwxmgP9LK6FA8Ln8solSTmHJg8+cWZy1m4V2yoZqdcCtrPVG/evJL2
vj7kLY5gixOphRJXny6WFNHUizfbKnw4ZhYmC/Jm1NKxPwaROtBnCI/QZACbrCWezCcycVaXLjuW
LoqevyBAd/UBMXIV//wRjkpooOF4gEjbJq4N+Hl+nqrew6rgfp2jaQqVz5FhNcwciWRI+6AbCpwy
HkriFop9zaR3LrOmW4hzCCWhc5ukI+uVpVTUCAVwwNtQffGCk6FHgG4EGoaufhOVu+wr6z/46OQy
U5KPu56yO0jy/iymzohm4oTfS9SzxJ/Dl2fyDSLkqRv2Uc+JxKnzmxqOtvt8u/Xgw/2xI6bX7Nkb
KWcpZ2FG3HNOP7/pCaMRsk52+sLUX/0gpWbiz2u5F8Nwcd51bJS/H2uvF2v6pDbhNvQN010q2bJl
bWsib7g5mkYih+b1e3R1FGDB/3qAwWs2STW+FbZa6xLK7xVhjzsISK3DUXoJn2lJPAnCkY+ZMgXd
KvoLr7IVIZGe9tGisvHMRhqOUuO1fgMrU1tBw0s7XE3aSpMfcGFxceCF2QMlsm6FS2t8UEa23uBf
Y4z9aV7ek9RKFxuKeQdFsP5anF6TWIwF3J0nr9l7Zhzu+q1tORJ9THiQF8K9NqlJryswfiRf/F0+
9bvMxUCbdDNwPG4BSIk9PLlZuCmqqMIUpy/mQPnzMD+5H1ydXXl49IM/OsTE9aA1JMgFtUu4CR9p
Vsbn/njDdEsnwM8DmNspXCEGu5G9KzDg0IsL5rqLY6ufIzcgam6fDjbl4YMMgyt7kkXdi/8w5ZzR
cWjJRrya0o+oFXGxO79Q6vfDj+sTQEDuDlHemvSEFOIN26uv4QO/n9Pwlo7W/BaTdJXQ9RhsQY2i
8W7ZUMzW7fkNpmXSgcv4v2vmCFmadYzipR2D2TnDCSitdQ7lrPZvAC1SRXE7yyzmXddJXn0lOIi5
8DinAwKOFcOnCJ5Yrw2fZHHOERM1ik8PjvMsogPH0/qFdB7lkMpdFNM4DP3iupF8TC3SvqQahW7q
veDAOTK4oH50lykaOFd/fm5WCom/Vt+f6mRICSycJfjTQGzBeYPxlsmbrskBHk1gXYnPF0EQqJBi
INmQQnhqUo+MbJHrhTa8enFudxFY5TUpMLEL8db5/AyA6Ut/xdgnUcneckiHE7RAV2qvA3UX63sV
t1dIhqVKyWO+H7YzsO7IwvdL9mGHK5Cl8wmsn80zVVCU3p16onAUXBVUsAHCv88MwuC64HufkAGB
sP06wjZAt2FerQh4HmpE572fmEnEQxbjyuunyla078LrbncfT9gpdT0ZXGor2PbIHfe10llCHcAh
xR1bwhxukin+XBgexCSXYaM7peXixuiWdk9zWGu21tZxWIWb/jQsxnHifzkF+eI7stFOnonQIECp
+O2P/DeTRXkzwB6UeFXHp604IpQih/31fxTysk+67roTvXgXu2JHT7xFmCK8apwXaUfdI+Frk3xy
QpMosLLLT3Ndf7w/6WTNh3B6/1s8u1qdCRFDH0WI4ncVTyjWz+aRjGytcjjWQSxu9Cj6O8bXq8Va
GaECrYBuXL95raX/j6/xEIK/cBuEVlIp+cPHt5CuE9C66dL5el2pNxFqzN4WpRz5/h/VRd+y4n/a
Im9h2MYs7evsWbu/lek6Gbn3zrvhd7umeUR1bOhO0B6wlhF0W98vZEa6+IRwiTxsvXdwI6m7lUGg
oBCXoolLnYOYh3yi+5cefA9IO5ICT5Dy5nqDuhCPnH06iN2v4xgT1btl89CEaLSBfpGg4VXPDboX
vAlt2u6e/hmWVI4vmquLWBAXTYHV5N9rJ+3YPLsRFWX8JGqH0WMQeu4AUv/ohabp5KhAN4CdLgpL
XwIdQzwZ9e7Oh68WMUjq8/CIGryms6Hw3uJzph/sSTZqJHZ2aPcX35jBfas7ORs3uvyRYHJT5i9h
wwroYN1Bvd1Iafq9KQjwH4xfw9JorLZzSXhvt7mulfuC9asGpvNPP7ZoyHfmtISavdIKEI6WQJ9s
S3OS94iKpxbPJSLvNHH7kYb/3S0QegnIA2h2U0AKg/0hTsjnpwcJwGCP1Pi1LbDUGEDhMw/FBBmx
eto8SMMAxmlUF4C2HJUdFJNnrL6wDAei1COTilRG+AlKkKnPFsqGnwOw+jpx10je3bOR4xXOun2Q
2xvkt/DJZi/HRRUlzVafArj/ZcYzzeA/BRKhJ9kQ7FultaUQfg0aAz3H8B+LiGtJJgVJatCkmbO7
WPR+j+haXFbAtwBublGhR17xu//3ln10bCUIwTNletfGcb484YWU3ZDR8anB7+kXdwRZl3TSY6w8
0pe2gGDOgQFtjJTyFsanolRm8hWmj2x5aqzzszPA5yTqVP4CnFFlEtR1GVUR3WN0rzsBcxP7DN+C
j4xxWE+gCfToDWDyReC/77CSgpRQcKSE8aPEPyDK2pRcPmJyQXRYwSYcuGxTLSSUVO5lZGn+A9nr
tnPos8kuUAwKDfxSY3WShJKWOzU9/KSNFbAUAhfjQ3rm9LKwLq+yNd1Ia4uONIrZYR067cfQLjIl
x8LOW2Ubr/WvXAyY9RrtvNw6cM5Cb2dDCC0kL6IdGowQ2yEMMygyHMrjCVnYQgzY413qMG0ChjoI
5h8safvKyNKD7DIejk0RxAgaNe9FVzXOS46vUcBt+5IQP9LDGAm2pGKv82oXGEoyZBDgXdNKEfAA
4Q5P+Ol2iaIHVITMeQWleEEeLakcZodk6JrDmwDn9n7ksNlP0LXUuFqcgq64UsvxBUYJlamK6aCX
LqyuqtfBV3LdN/y20Bix14Z+0ZnnNH9WCsTQ8UiZgKK2ShHvrRa3qK7goKHs1sNRt0gMPGi6aaEB
gqFaDqF6MB50p+HC3im4o3qs+NBSLiaiOeezhsr1KS7zM72FWHNqSQK8vZX7r+gigadJYYTIB0QN
fXJxbspqUctcBHNopKNbf2sb4Ut+lUmH0XHJclRLDC8G3U5DWcnlGrsZuT8CdAgwIIn3sXZAl1f2
Xku4+SMdI+g3B0oPKPRqeoxffIrWZGiH+fbGQGWs3jT0ifOQhVGdDcYWL8pCMWd2GGxLoIHtEb5t
yIdL8oGjCqvbIVobTzT7LRAJFJyvSC2LeY9anu5vofGcvQ2MK4FVval3ok0i1tFKCJKve9x5RR0R
ZWTqXPG1OQRaCihH0PA45Yp5M4ihEKBMGNV8y+w+495eNFhDswg2bbyukar8InZ991639a8Vam7j
UEc8hW0jPeMCsbtVmIuk4fArgDSIDbYgBU1p3drf+RR3WrZijyXGnsjSrpmddfPBXsWJ88fBJjub
LVEIlK70NPPIOPRMVD6X3onF5JDj7g18XSnNxDfz0U3dyLTSqRQN2l9e+B9pX9sPsTq1Zl+tl9LD
+uh59aoQ8uMyP80xDIbvfJxfmSjZ0Ga67oXalZyx9/dmObVbwrqPBETZCyQAA3VHVYVzpi4eGC2g
clpBrtkW100oAFneKdclh2uEFj2JOii7L2f7LIsw5Tx4CsuK0V5rirV26lV3aGUTebQazkN0uc8V
w6wHtqM1vER+cIj30IcNm0ei47QHiME9zyFU+gmeHhMgERrnzTEFrkEVAbVD/WyW0WMBLEdELAhE
IzSl5oOauNXnauuI8LGqWxl03rxnPb2esOcMBjG4q63ma5De8xZg95q0XgTILX+9AVlGO6+17gEk
rcl+q6DVNsR2AlmIoGYEX7ZFTCX8Yth8NeR+GkHZDHQ6JS7ca/1hkHdRWUHIknsBnSauenZUkPjo
A0HS2UgUqVoT9x84+oaBsn1HPdcParXOSkyKeQU8ZpGIIGzE2ygo61RwWPByUSlZBKz8Y001vX9R
oObj4z1gGPjoadn2SY9Kz7JSLQcxUGNqHsKN3km038jawloFe4+aaHd2m3q1cxZIO1q1GLW2+FvP
56u3If5ncFC0QagsSAMzrxJC4Deor6muu4GzoCczjsFN9V1f4VdIRLxotxEpRYzv1pfWNOeuK7Db
Uz1IJyFxC2DSyCl2rm+SJHj9bvk6+7/CwZJRISTY4iQfkbW196OrGRwbfkS1JdHnUM7NOcoI+Qbm
GIGoxtgalXaLe8gyqKDZL3bvkEbOl/SoUX6/A/aKoSidDsf9yAqGCv9SVlkxLplREyAaOvtWiVHS
i2m+gYuCTN5r6DSIs05cE73X25Ov+Z1f1O5U9f/DxyInY+4HiMcttHUl/DqPXIx6MmhjSrRNOLeX
cSq9Z/3IYfMZZ1r/3ziYLfVQtY1sQxAchqxZ3gUs/cINL99PtOZ/mhWxp6dP7zZFYVXkqHMaEfZ+
xycHRPMq1zxTOuZo2mvBWEd3nnEKnsY6uEaEQ6QVehfYYXQpQErYDt5qO7i/fo2wWfu3oEZajd/t
eSNRJK6WfjQE2yAtagGh2oGfKWMijxj4Blmy+qq38pOQnjrZZ0oZPEknTFCEMhRlxW/hn9EaXmAF
D8IIPTwMdutq4R1vajWttx8klSIzgiTfp0Gd7vlSX5F4HtRYtApbIgvZuH2gN8tgbvEppHRC3Od9
wOk9TwvyjrwaZlUdYL0aDRcFOZ6CtqIj+ycEGGcNc3lICNEd1ZqStgSvA5I4c9p2+MA0reniHXlQ
75kYW4lJX9Fe77XLz3CdU9zASe9R8WzWUqJbhkYjFQHD8dzMBT1AKR9Kk6kNn7oFwAHW+jjj3CcL
H6MtbKVAF4G1uwP7NE941pm6y9/qjyfw1HPGfY4ZFpKbpptT95sUBMC5UxaXUJU4lg/PnfjDT85i
wZy2Qn8sRHTrFMPek/MdMCimECKN5wJ6uCYxPGVd5WGAudX3Mie21pbrcDvl18Y2dkWE77WXWasB
LjXoW1qdpTEryCfQ/O+insuqcxrs2zt+/d7poSV2rp81W8zfzfwPWw6nFFxu2mOLqUVVO1GNjYWC
udljJ4nXy/uVLNuymlvBvxcI15g+Hl5zL6iBAfz5bSXIGW+6M+85qlRVtwQFM/yZ30CJHWut3kgA
loDdwxsziwo+5AueQu9DjahQB/8Te5qq+g+IsnIOxpuTJuewHTfwUQd+3VKoy+zUe3bLlxnnUHfy
WYzuMFcAuQ2mdg23FYB9d0Wz+U5i0F5VPoCwA5py+1RujpX4NuWYMRossY1rF4ALb18HqhBcOyyD
VfWiWLESvsTZQe/zBhjzrSeu+npe5l7nBAzfHpMxitgckdf7+LAR2BUxn7hnBApEeMJjca5Inj8w
e/fFpVICdHk4FtpHuG/hFF3eVuP94bD3bDc+s3BN8i7hbMFZSJUEbHD/78E/p1tMll9gX6nHOfBp
L1Gz88/G77CHiGCdeYhC+g5njOUwVdYMJ8Pjdm9vr82XEzYZoIum+6CeMO9O2xg78R/+dyF7Xh+l
aKn3W/8RUyri6GniuzIoTni3prDDi0cysvTCzyWJPgqcVcDWHqfVNM4wbw/WbuTNH7aRdin+XWfd
TbyZo4BWv1awcgoT7DsSSo6KDT7VKBkXuCHGloybbMtBOipYn7xT9zUw9N2vZNSp7kxAQWhJ8ZLm
PstjwkKUgAxTLjOA0vlR1AYV+18GIswITm5qwyfIzWtZ9QYDSaIoJvzdVWIouwy9a5aO6Qh1aRnr
J9pl5ZnIlCm6y3hsjSCem98Uscp2mFaS20SStIMzKVTKiqDySZwbaQAFJPdkg1vepFbKrOc+IsnJ
6zZ4Is8JZZixKwC0tAn6mR8OHZEj/dnqvXT6yb3tzh+g63c3K/AkhFl/abDeO1TpU8n25hzv/5E0
Pp5bok+E//VkoWYUiyWFQ8580CBeH+XN6IVq1I7e2l9n4Nap/BXXgtvPrxili6PjZxgMd9voXiuo
fTbfH1juZ0pZXhw7aytwso3DP1JHw3tuGE/TxaoC9I7qwwkDkcXh2ptJzX8sPaoJ2ROGkTvl2wQB
cWLPlb31MRNWc4Qm7xaDji/8gxSHUb7s6XjaiJBtFgIQDjPa62dJFt+6gZwWn0Q4jc7e2006grH1
J39wdZwSYYglDpxtfAlDBQmHN31ovwhmYu5KLIGHo+2VA/SeAXuv45A2y9Not26ZjHp5L3gAZ6Gv
akrrn1e+rkjeVgenpAoaDjYaHGxQdRYhJzlmZl5XNMfUgBuZFb4V5ecxKnBembrbzvT6UJWG6ji4
Y+GKpuraTbxsmp6swI0FFEApHoSf6IazFKy5IWTwRQmu5VBuIcSfljDg1oCBm1EPjkwawGCHv3gd
5pL9NFAOF659v3zdMwXOLshKVOOWQWERX/V31DwWlg9RK9TrBpNe8tCQDFCy3iyuWIyZfyJ0HTqR
nDnpBxQWlaWMDf/4ENiF/6s2kUMWeIpwBBH7+XgdskICqYPaT/1us4LIsdob+j1HbRJaZsWUUH1I
y9Vs2XA5OmEGqQBJ/Ajl5v5gCo7v6Q0K5WJadkRjqkXdvACKpTNuzwt2Vhgp2f8f6UZpWh8cYmKK
Qo6mPY2u96drSgVNKp9sxjrvyH+NAZ9+Vi6yKuJejaJE4PAUfN/Qt7OFsEN/x6jOgRYtlqoZJR0Q
8yzhQ2gpgTp8ALouoFUp2u7ZmfIBGKjnqMvk1XJyfxvPcW3Qq7rVdMZE/uS2RLVnXK0zelZTzqbl
bt0yD1S4Y+CGnvQsMIkpy0SSkTt/MjBbGxbG7m4zeRsemfWTW93+BjTdM7Yb1MvIY2IOpx3rQg0z
/KMXRT+fYBJriEmStEwlwFiOJHXt/7nHX4BgDCt9Gaq4iqun6DKlElthMQuKAm0Eha+UzpWZbOQl
HabQs0Yr7C282fhBEbx8f1oY6Nb1wqJw3RXy+FjiXcujXIL8+jZ38A/w4b2lxvVVORF2atlvINi5
y8EsKOdpMjYTuaCOrJEwM6TFrR5E7qVIe8/EoWVOMnFcxOcRjW87sbQmGQ9xH004nkWxs9/6Pc/J
MQbLSW4wxIO7b4BII8cDGi6r94uEOYZdk8gv1I99WJx385g1wafz9+stInACTIRvyX0q+ulhg3yK
HBEuTDiuRNCIa4Z5gpH/B/a+Xn1qBvr9TIUBsoWwytSg4E4DvTd98J6ktQes45Atc8PcBJZdMDF4
GUN0jt6JnSWUJTCq+FKIwkPdI3VGRQjXseN07NErNYcWKP9jBL82vZ83oh+Ixx0diJPSFQ/enMp2
aEujNhprImfKusjan3K8YjsJ+1Chvv5saaKk1BBiPyxrN3Kt5oqDOKjpeRlxW2brv/SmX3v2LAfa
JWsty8kXfKqrOfuSAPSweNxnhwCU8zYtNmFmYnPvhlHZgdPtqT7f+/BT+Y9Uwsz1nFY+hh6R9gfj
TaGxSlU3/qrd9ml+TZ6ffyEDLTrTT8fAC/241Iq2hMXoaZFzeMl2QwpcZIYdW+MZQLjSph96ZEfa
4OHnzFimpEEWQJelkFgLT7eQ2UEfiFDzG2GKl6npKmT4dd6RMTPYDpU242G/OoX2DK8SKzZ2yHLc
W6HVlKYLkV0djoNypfc3dmM7jh5oIrnaleno8dOp2zQTOfpg2UerikX3FD0fK7Emf3zo26OtKNUY
4rahK0/bjQ39XaXYxhISHt6qBy40U/KXoGkXi4ouc5LlUWzzZOOd3TR/tl1yNsGWVeaJ0gyYvUou
XZZM7C1kJI35joVjmW2tJFaTlNTnW+NxseS1pCodx+LXuB9+RYXE5c/iIMfR7nvdVZZaAg42LxPg
izAQB9UTfDF/Rsy/t1yLr96eriGDwEwsW+1DUMpN2tjGrzDuhtujbgUIBi7EUXdd0wz8L0NHffL5
qL10EDPvxkCRZtdPsM81Q7xYE/5cIph+2vSQ3Rxs8GYA7HpXF/iiapU81YIKdHLesoVDkWBsSGEO
EVPMT7fOYEjasIIOqNEdbxMvsGFooB93D/22xuvMRoeSZ/tf0TwYxdyLaR10i9IRrbpGxCiuVW2N
H78xZzhUV96tWUcs8MZmyjudSEdbzaIXE0j7qTldqRlg6e+XRKR9PeDIqXxXxEuP1DqkNlIZ+XPZ
5wrKXl1/DtdOHp8B+A90XxA5uLqywSI17zEWaHFQotLUBBVHaOBMLWPkyWC+Ua9Q1/Kt+KjOr/zj
tpsOOXIBca1I+vhQs6bX7Rh/WNoCv9xEuIP9qCc/YaE2Z0K6oaO4xFR25djinWKEZ6HrICf1mkI1
l7AA/a76X2NFPIlJMIJw1hiOgjaQT6+vg+tZDeIP2CZKFMyMxXqDBSitw0LEVJol3acFqW8M0HTC
tqLYSmoNu6/J/qd87FEUts3tJJeitUTIc21YikjdQiUhnve4UF4vIgy8uvcYoQiVCDlha1dh2Rn8
f8VngDaSG8GgSknp2aomxt3AQQb+4hDXZwyKhcPvHS3z160h2QvP8h83QgGNlTvlgwBaTJXZ4kW4
I/OOTBfL17GxSgk5z4SVqMd7npn6dP4wMKqsOvKCOFq6yQlL7bW1lQx5jKs2QheP7DQqcH0dZrh0
wCPOx+M0oiIhu8qgOx24cnjjFNiB1sJJ1Py9MKoybqi5aICpHTKt6VB8qXtRDMN7l2XPI+ZJA7A8
2T0rb2UuEjBJi27yHDfCc9M7n0dBk5JwDQtECy6enHIOQpHLq5uQIsSp//CyllU8ZNs5USYJvmUg
P/j7jC/dfObKS3vaBeBpfcf2R7PuXlrRaeXpU6fYgINzYBOrzoizVK7qO2697qXKP+mQxmNAlt5i
Jtw5u8LXLvnFUu5pilxjCRaNQvMnM2TGFGKulgcmBvzaEl/iiNFhk2/HtO6PVmwbrP0NugYN8lJO
wWLm4eU+Qvdt4nJs86GlbNg1g69NLZQbvPvv8eD4TTTNOmYTSRjYl+rdMj102f0NMa1dtSEOMWPt
dG9FTY3v6P4D8cPcidFVt9R/KPatkGEfZMNcIDj7A92Ip1W50u6YAF0+EXZFm+8H1KWslX+MHsqV
o/cc+zKiunsXR3+S1UZ3sc2A4xTunZkiv/1YJHqZ8hwZAgk3wflprSRurxPRFgYeDVXVwRiBOC40
iZg6bkDQJidZ0PfYNcr6LykidPOhJ+dO+DjQ5WQ2SXLj5HbKy1afgi3Lrrn66YL2pbX+xpoB8+yN
RCsOpb+ip/2rLZl5OZmeJP5Ua4xljjfeFX59s4lH35R9fHVFHCGzQHvuZ6RQwH83phmBFQq2WX+c
5AxbSaUs3f5euf0fPCOzm94q+/VMLQZ2F8+TvHjwy+JxdrHe9m8mAhIpKbpp7fFJS71ZhWE5kcp9
SI5bt3rMJGcerbC2UsgIcLYfcyz4ocWUgaHvc+ScDI4loVe+q92u2J4qWhRIfzjBy+k9vv7hDZbo
CEufbpB+MCkypQPd+wX/p67R6G9xeVwo3YxxpkuwrNlOVK2hxFly68NUWFdL4HbgRgsWLkd+KYCf
UYQhPq4NFOFbz3bePb/mNT3tb9CdDsU6jIY8tqxAUwmnNmXqzUnJXISgNQ5DBV0uFDTsvJ9As4Oo
MRrGhP20YMY4eDGpg4TplMAoVGkV5BFhQWdScq40GjMlRBp809HAx/N6FGrKgS7lhqtvOTt+e9XH
HtI1L2tlJl2U0odE3CitvZCDmCS9R0Om2ywFqIJJoyi+e3+yg4YR2UCT14J6feYCEnkHGO3XPQsh
b72FqUawJy3gPw/W09XgY6yVT2EghxekOuvh61x07j4t0SFrrBJ4lBGIui8NsVjTJcO9ycgs/y+U
8D5BuIZtpC9cZ+jrGmc+FV1UcL0YIC3v1rQ0z4VGRcnb1RTvdS9dU5T2UcioH0NFz/5zbhhODYq4
YIlPgpdXcnuZedEOMIE8hQCf3KH02EyJ/YFhOPfJW1afGOlJR6O5BOmc+JYCPODDdSIk9bMIPTVE
kIcyHK1ShpJEXqzSJRDVyx2KGr2dbiCePC9ZZMzILBBZd/Os7kTDxn2z2Zu6TqSJ2kDxnPho62Cw
0KS57ylZWeT+QM4Wj60n8vmoaUfAmpCsmF435x3IMfN451DUcPPBNbxPpdt3VsgmvJyrIP/ZH0H1
iArCQMCU5VupqYCgq433quPxPhPrjt9HL1hDucmQbN7TcpySi3QE4BV2s0ZSxCSmqIMowtcctngf
cwanT6jUpk3b/ihvLZWP+2mtMjjqDt5GK3X/VK6CMPbaN8G8kiRBPyT3Hjbt0tqsaeo73YUmWWEl
bCanmn9MUCbH7xD8TWiQmyAjYnbM62vNci43sPoZ1JyaNUcoi4vIbp52hN/n6O3OLj71AilFlR+7
zGouRW3AlLaUNT/ilNy2JPfhpApxsZeI5ieZRvadLsf/wTgmENKmR6p7ayNKKWUU2kLAWjymOmKp
dl80iUWHVpZ9WwSWTDxagA7ZzBi0lIV2nwNk27SK4b2x8y+rtTOWfQhQtu30Crr/VNUOtHaRNE0P
rz22H2ol9c1l6tFY7PxJTxyXhuARdi0ukRD2ARJlnUXFlpJP7a95Wc3Afazb0q5UT+1nOwwBzHLH
Z/Y+s6uxUOqeXPf46F6RxIGMsH6t8BqVhm51PHbXwLMuuHBgkAXqt+bbvEHZgCao69UTsrCY8/7z
5JuqAkDB6rz50BTJd3mLNEWIWo2zuFo+KYp2DuvPnHmPwyTG3PN2CqXFUZ7Q5ebphOTVBFO0CpuH
YQub4nSlqvV3POt5vH6x/riSVbCURbXm88lJfCp7yPsc/AqD76WmlPa7/LF1CKIL8RD7L1GzOTRc
hhMQoZ4VNPac5AXDs+M4QvLfm7IFVQfoPhP+3kkbn4zx1Ypm77rV/TAf78RMIUGzrkVYtJtjtqEC
NUzqY3ynhvNk3CgKntcX0j12DfCVA7T0gOj9ZSXpaCobFNXzy/UoNPAzAwHg3D9i9VOHVG2S5e5E
aPHWyiBApL/oVvipVKxt0RbK31co1GLpvU6cVWb2zZMUU1jk6oaixDFStEXOv2kXIwzSQZjSBleN
fFHTOcZ9lAv7mXR1ipcwBtX0jBrPVZZhC9cCvxzWwESJlBIKwK9NzETBF4Nfv8pCc6tomF6BDiNX
t1cZrnosvzMQyjhuhfNByczXaoJNgYgeTzX6UbzQ9CPc/Zsrz6p4ZqRWwUWI/8tCqCvw3rrINkv9
uQuf11gZ3YzniK2z8wJVIk+xmmgPujhdRQ2byzdh7twU4MzKbUqbSqHr+i9W+eE0C5d3URT6ri2w
PVR9RGIQKxSB323sFaSFlui3Tr6/EUNzdeyoyJZTXxvBuO2Cw9pqLRzQJ490zXW682W6dR6S1H7s
NTc6feiV5vHt8+CRDuZwMt7I656tWEyG8uFqAzCoKut2aShceTKSleGQGZ+PT8+RJeJbjS3QhAcm
yeMFUoVbbNA7EPotByIVGY7RGpDnkl/DgtukA11fQOPyjXQe+U5UVDUavDo+k4fyE/cv+B8ZhQ29
g9BL//CMJHvqdVcGFE6kAupOLduuHQv7YYtOKBjH6XPKARgDe13tnW80v6oqMY6F1+zerYTyV4wW
dX1I4MnMEHhWrOpYwmWiRhZRSXPN1oP7pKhY2s8hnWHrRorD/eCV5JLvCLXa6FZB/9ozb+HiGrJx
xk8vNhGggXIEN87mBy8ox7RkzPzlUnyIlD4tSkiQ/1DSpORgZiZ0iI9a24xOuvRzjFy7ASimv8Ow
G0W+a7oKhqKnx1efE52Z7We7HOAY2wbEVkcLI3y1b35TQQvX0f9sQ6OcXl/TwmpseoW7Up06MNcg
UY9tHHj5j7Tpo9yTO7dZo42i31Cx+2/bdPxkEleVzSt25kbI8S/AflSlzgONmtXLDldiQRLiPDrj
0WdVwD0IfXqRuPqIz9RI8/VSfpm+54lAu4l0xuKIEOpxsol6aLzmc/jl25NguRg94leprIeXIejV
SVJz6v/kjEza48A9VEpAvQJUFCvetsbjJAVfrk8Y/oMHZrz2cdoeIesyP9OX/pIOMOzGeQ6AtkFn
hd0hmtKWZmXe4TBsuIS6QtMrDsX1JhcnFZq6SQnSY9zD2p0wm9HlTm4utE/gNvbM9NuyvuHoBAp9
3HCQA5lnOFmCN0iE+DY3YqzVD0UuDZmcbaJqCBmBEliQqZn03O5dcJwLW4zzFslYnk0Gg8Yz/q+x
7NqtlzHFG4i4cGrrxOeIsVBWY6vxZzUWSetY7UH3hnXou6Ao60VjA2US25UVuIH0exUiTr30zrCI
nQMDdtahKEEV85MgCBiwztHLX3owvMaHu3nmzleJpRNWUv+Kt4LyXBl1QEfh4R0TMWeifgodRvvw
TOtykOYT6XC7FbHzfFf9dc2uaa59P+l08U/ZfauyCyvQ7qJNLg9zr1K789Wym62y1yYrqlj5ZTM4
znTs/Oeuw+L1ovdGxuZ0DPIRsju9I5vLP539dw9qfPmLO+sxAslIA/X+ec0CripKeQXubBGWj+pm
wJwNyqFRTdkgIteHUn8x43dNqXy49D/8cBCXq9wzYMDs7DGqEpurg1YyJaSPgptg3/nFm+vNKlmD
x5I7davZmom/4uKvcXBkcANrX0NIIZVb7Fkp/AfyIJoPFQTqY9MQmLoyBNXG/b2vkQpwRdn1AC5I
UWJWHXE0tkn0RYvpC08nw+mumnxz583/GTM0OHy/a9bnsn/UwTpOxVADd2FElvBO/uniXEOOrBZQ
SFHJVak6xT03AwhV/cCeAiiaQwRS2noInA5jNDmpEp5nBINxxy9g99sRmortZsQeJABtwVyKJG2V
vryPpIoUTqWye7/pJoFvoYC59U6AFrMs1gMVbYza1NQSmqjAdGhrK6EIbsFi1t4sF6ZhdIUsqOva
pUkDCrahbAimdoT1KnPaSvSM1Z5m9U7/hp7fSC0kxGO/B6h3aQsDq/Gi2EitBFaPwdHSvVhyC3Nw
McOgyU2SYrJLw1G3uKhDPqZXE3vDZiL7ixsh0UHxFY+d8bQbt3DY5PjNZ7fPZYEtK6HTR7aaprwB
evhCBoPbKW6KAzJoUMweRDSCbf66sqeJjhCY6YZ0MkRvg7iAf8DtFyzD1p5q+zrA9wO7GOHia236
TxA8z2twZ0Ow0pZNpEgUE1ggDBHO6k8PLmnSBaRO1ReFEkKU4fi4OV26+l446iJJzN+4Z/vysfTM
zvBME01tz+je3gEzKiM59nQJsXqOmSfOViu8t83GLWwdR6bVBPm4ZIgtZMW4KAcKB00wNjoMs5nF
z8irZE5/Y/l2sFNH+nEj2mqNZyySsmoUM6+t8dTZIRB3xwUSv4BtO77aN2i1RpYKSi5phO7wuzzk
A261FuId8tbEyHFY8r/lB3ymoZttLKc2uQhnC/V10fBmDTKDw7QtUgVYHnW2yMTAnXvBBc3nNqHE
egnBWkjmhRYqEdmUBT0HctUfX9iPJGL2btVIih6tOhkyqng6qe1LO/gLB38Ld3u/RdDYtpVauQDG
kW0YSpqLM7ut9NMyznBfUcIPFQ2LT5fnvc5qMzIC3gi9at14dfTTL0dan2f+m6KM2/gq9WTWFoTK
Th1ZTK/EmRLAPvPaUMEMg3/8H0fwTPosvecFCYkf16vCZwtGxbYJAwSJuS/ABpfyrrUJlRbOMh2N
bdBuHA5kw/+NKEpkc9+KBZwnoaT/1TF65TL4+MZAP/HrOGhU2h7De2gehIB1jgKUdSa5dJg0Ae3K
ZSEG6yommsGM6tJuCBQnwimH3M8O0bKn1/L+mvnotChXWRgYzSEByWvIQLj9EUPFdHYC7MEYyQgy
4Whi2rncv4poRtg3Oas0C+wBDGaT2nRe/SjUIvgUWrAtGLdBc8swdjGAHR7aA82MRxx/s8XZ+Ndp
2htUnecJhmh4w/36aPgMXJfUS29YIvg7YBBuQvAhlzARHT/J0Hh7i2yqaA0RHqnL9O4qzolqJk4o
m2Ju9SyW+ME7sC4ftyTHwwLX+zwpASGy6Y4Z7ZmS+P49IwcMVW6HTM1/Ae3ak/wmR2Onrq+Qw6zj
ortJiCSITQ/gI9kWnfTBR8upFqoAXlfOGophM+SFfq+nR3YSaergJOr4kg4zRG18srPqmxBifXsx
MmGJg61ma3+H85oQeDMzJfTSMGc5aF+DTISLB9D7QEW5+RCHGttW36S8VS+4hOVuhRjd/Ni0/+R8
i2qlfec+GIqQvZUQEcF4HgkLfQasM9XD7oXP+ZKcnh8wq+wEOIj0swt5JBNzSV+s2JOaw3Jk+ne8
JtqIOIgTpKjCV6SPa5nY5+xPG5QJ2qmiJ38bqqv0dKMGK+6ekB/3S5RBB2gshDFAS73F3pFkusVj
yM1VnrBTjqLh2jfkzI0RGTGf/bH17BtyeXmuF1Mgz9ETDVFTEDlamxh1ngB7PLuyH+i22UXiAaqC
T3Mlt8jb0PAn5KknbNDC3z+xOeg3zof8ZjD73B6dizPR4IOCn8R9/nNHrxkMDImVOM4HKZSbkwuf
KJ24cQ+Dson85uek5Fz2kv+lAdXYs5c9/9ChT8u5M+ei8oVpY6OgCRIulQrCcNoBr7F50P0mwNAr
f7N3Ca1Oe+cxKIMZKdXucOixKDjdX2yg9KZaPaUEIcBFQ0BoDs8nsiI2vEVlmbP6y+1YEoAOcvxy
BEk+wCPSSfdIemjBLPrfg+SFmM61wJzAKhWo7vJeSiuzBzes9HyhhqPZlcpobkmMZYGwIbBg/a3q
CCi1hJoKyf3wQOWwwd7sMqV8yP8nR9bq5nsWmX9AjHQNBpNv04SS1MSXp0qguaSv6R3qdPp8MyVJ
I1owzK4EcY0Z7eT8VVwd9fZUEVGTpEalvPnc3MxL2yc0M1l22MuqAffjNEFJxm4I7/cqG2inRtKT
oscWguOO+SuxO5wKzJ1iTmKlmrHRjTPtf4Xn1t0F08Jodvmd8Q6jRGsJSk4vCJWGwvhzttn6MUFi
zjzG/bc1Y41tHzXJqfi20wPKsLIFCnkkKIOxo36akNuL0wMALHNjgKauvCSgfJUV7Si+l9zIcPb6
wgugmtUHKxlGzgLBrVSfioq55f7S8A4+ubuSnBjhZQrUCo6UjUufg243r62l1N9H6RArI2wilhNs
3EVVHWA4MFpTGVIsp19bSEgwB5+cXzvKjOEJUN4QiF6vzyeEnv4dqkVzyk2gFD3I4bMCTTtYGISg
omKIM77dw0jWELeRjnfL8njrAqkFLkUZ8DkiZ1A+18OBF50LsNhHxH4vtuv89sF4n11MnhxOc3wz
DjVQIlSbpGaGAycBhKFEuXMkbu2uW9MaEx4hO3OHD87Y/YntncoEQCVebQZhycs89zb7UVBbPmI/
lEBjR1W5ivp4NlrCoOeJed7jzkElJ7/LTKE0RS51d+cjNsyQD9GRIzWNlsKSGJZp20blYnuyxMQ2
It1xvdICh37jSSaEHa/02nsRB+Uy8xpldxYQ/yGjF3T+4BvmwbJbM799KFU9PfJCtme0v9JknSi2
gY/3nkiiVuzxooSipBTObWyVwfNwKiANOXVM3xQEueTKSkro3bjxQ8WrpXJpFGEKHk05nJeoOHPt
/DHLcI+BwWwhI5mvcR7WlJGNcIIb4X55gPODMP8OmHSMAq8Es7IGOwZvF3FESRG35+XXDXDQ1xAJ
RATxKLj3UsJ6Ab08gMhiySE7APHN/lRyUDpLLHLBLmQLdFNepD33w2TesUsvu7vZ/8HYUUww4HN6
/4OYP2IFHoVyvd8c8fttzpezre8BMzECWrKHDqBpP/8FgJmjeclS5Ap852/tcmehQBJnqEJgy7Vk
CaWmpyyhM9QfdDrvIkAknxpaG9dzO0H4Dvbyw3b+MPF3jg4FyLuR7hJMt2mB/CtX8nxvqgLqtmDz
AmEfit0EuZUbruHQiC3O7XSu2ZoSBVt5rr0W5zJzhpog8EYu86rz2atCailh1YV6YqiPKi01fLGW
8Vzzs7NJw/cSzrpUgR3XrXkzEmQNwOBwV9jK1GT4rkraCq2Lo8NsaSqqx6QV2a9vYsf3aNYrTM1d
Z66BkFnAWcq3eT1M0c1ZK9Oy3CmFp2tnhJhCuuSPTKwEKTs+evNdsxjiiONYp9pfBGI7jATCexHO
JqrYE5DhAxr81f/dOypyCVyy6n8jonIbyGr70XYnyu/1Rk2FeacIncPd26sqHNb/Lwq6pYfw88Kk
dz1z8flNFOSruhGLRHNy5+/9Ewxzgh30z7jEbtNUcRZ+GicmNBXxQYuZBQ+823rqNyAoA/Jiqjzj
ilv+JYxCgNzRjH8xgS0L4Mp6HjAuVMiVLAkjWZzu/7pRerJ4dgr2HfCF/AYwlqHc1xCBzvmW8kof
xjbjTvDrjk2o+BU2xDsf+Kx8CcLvdz4ZaGHeyviOaW+3Kqupo1fPVaiZWsY/xMC6b06B5iH0NxTG
1Ph7gj+2AujZyoUJpCt5rfySVnkJvuuDc5fAG2KT0sl3UYHC4Zr9Wf4+91Ne8UvHOpdryjWBlzSe
ue8mPVm2XRkRaNhctTHtRAiv4ZclnK2f1rBi/kWZz563hRJZfd4OEKyggGrcPaxRxSKXq+kHMhq9
603ikVjgJlvklipklXVhilUZm4IubB/sNCR8Z8oN490XukWU77USM8631U77uA1clRP4urajev4V
EWFNxKegE7jPfazBimqqAOz6/mYWRYftCDbA0KP/g5ZGLBUKnOBj593+iwNJvJ30Wne51fezp+Wn
6+WT7p8zXU3EmrBAQJ2aX12iyLSlZcnAjMr3M68JeLnIcRFYO273mkGg64AjxHWfqrwWqeRouQ4C
lahAS9LSHr8XsJR4OojQq3VlyZErNCDo6utVk1u2/EI7gKYcz/r8+Rzd6tsgOvEuVkRygxV7qG+2
/U+F/TLp+QDdFLsGVxJhWHx1o8FhYMv1gjs+lUQdiO1PLc9653a0xrJl2z8yDVV/UT/kM7Cgiplj
lizpnKM/EnHbWGWok2wdky3/wzwOctqr4EApL8Vmu849PSPysXa21mnOINxBAvcTUseH3jmWHRMe
Dc9AcUkQysd1Vx0s2M6g0+v6W0aj8p5esuUrah3UkZ0wPjW7qvm+ucVv6yoJDBbNyzFEDVsrEb8N
ABGPvpESYDeLp9ssd30STmS0lDnnJXUNXvXLe1nfFjgTX0+6hzV8EpKXegBc/ZJ+0RoOX5Oc3mC7
//wAIGrEljPAUI1TLjkqhc4vHQwfvzGeCmRNVFbBvAWKFpLQkZ/p4JD0AfapKci02t8gew0hDmr/
NWWLos6VOpDS3ckqCcRtLYjbQSNbDgHlArV9c7VWXXnJFONdb9ujLumbxjqleEDplHzCJjRuhgRq
RwJjJhC1N9g+GHGDH+3wgdHhX9VXvldNUub/oqk+ol25NQaukgOhmQIBN90E1CdZNw+/aa7aeTyT
Zht8oxdPBRI1TYDn0+cYqcPDsg2uKdynKnHG9AXVrNQWB+TmpQEj0uYIQtzgwfxwvu9yvN6J6O4f
evwMZfQF2HWSd/RC+DG6mfjwHiJcFlgI6HhR2SVZpz1b0EMZZquNPZ2nCx6cTvTEkq84PYzzDD6l
DjxPCL6HIs9ROkrK1k6NgsCmIJVw2PW6Qpc9K6VC1fscdOpfL5QdMRQG7K5c7zx71hrW/tvZfo4z
q4TLErRyofWNIll8V0T7Wodc4FIBWPQRYSKGSkTX5f9HiWIioJTZ+O9gtTGYHTliRq4uMOYZmQVU
LKD6t6MebqWxImPP6GQ7o1wh7L8ILqyY/hvWG/NWetDoyLR459xs+qOjOn8zlYsIqoD2LmlbFtdQ
cMPA5n1SlHlFiLTC4vuR1Ni9axckTclF6T5Bmm8HhdrjA1F44HlIsGVNupgRf30n1ZWTrcmOsL3e
kSQZkaDv6zNIu42hzbHO1oLHsvo7a6xi4RY93gXBm9ZH10dP/8RyQ+9hJLRwKapjSA5QklI1REH9
3ksEPNOzYRbUmiaY3z6imtioAUeiEHf9hreoU5bX7/Hlg5/5qvz0K8oRbunHNLzsmaoq1ozmwZu2
Xk0DIoAPUa6bpSPD1gDGMFGbeJgUqtk7v2wiO3+kCk3SIJTqtgiM1w2E258oor63UsXzKLJvmhga
Q53otRIAaNzinNCNC9hXWGeUTs1ObHrr0RcgKXxhC2O2ZBvd7KVAg8L/29F1PH2fnrgF9ld9zxi0
3fAGd2+U1U/J5rhgs3ta/xqu49W1Imulv/5xEKN3RMTh2B0lPNUBEZolaXynlDID4FIzLlOQTE2b
wXAMJzBh9Op2eON4+imlHsgXkytStSSOnQA82pODBux71Q3gRBGXn5rLgrejmAJpnBEdLbiEzVHx
TKp2txtbeyJ+QPzL3XDVAosXRPwi1hIxCOTKc7BrURqwpxTNb7WktAdb8mI5/ibx6L1RBBoLEGb7
ktPX5cOjBvs8NceFRv/unsaOLDsAqkleEwfNdo1Dm4jqoeF+3H88nQttDwrYrKen1UEG+ityq5bO
bF2z04D2GuRZNTg0ynxQhU3iPPTC1LF6c9jlneAkvXALP1WEpN5EsVIMVb9lpN02JdCyzo4tx316
mjWM5b1Uu5xlluFOslZwx42sUnbjL9bbib6E2/wyYekB2VYsbjqXdKWuRqNYdxn14ANiLBquJ1b8
xVS5OXAFAs9Bvki4qzUPRDbuXUT/1YfZtd/avuTpW8454+1i5Yycava3CY//Avjd6Nyh26HGKUMf
7e7D6WECeXVPa+LblgOCJLKVPpENinM1oCC+oPn3vozEsDPw2lnQpa12Rct3KGyPC5f9I386oq4y
wRGXW1LhoOnMCgZWNZcZiQIqux2V+dUTuFBNQU7PSYWoGz/kv3PVt1PF1/I0ksnYl7+IIb6OerZ1
3pykcaorF9dORhDUUoY+mb50kGqg9n6NkY6u/+Z7vST9cyfxDuHcLQBdEsWeGxcaMrc8mi4YrAnd
mtUmb3/Hwf7flJRqaZOLC5Nal3Q+euBymKWsk4zhevcegGd5HKIH+jVDIVcRFuYCZd563uWXD4u8
YkzA86tsrBhI5qjJAOzs7mkzD2UOjqdjnh+eGqXmv1si4TaLvP3TYt+UYUyhbLFTiSoB/8igJUDU
P8W6/2m1FO7Tp07gRTJ9AQNGcLQrqsbup/YoztzB5j6zJAT2MWw6fwB9C5eYPQLlSKGV70ht8Sq2
bkUzINOerXSPXxyMNDbbPCQ8auljNJEDhSLTn4X0D+qPzZcWC8CwHVH0ixD/jaB6Dpgf1ViGgro+
tWRLBQagA5p+e90pr5DD7LL9RvlVnXZpoxNaRmPdihnhEEiTtIvKRZ/Av/Y+viZ4UmBuLiTCaYKj
mBaRajouBdOPGYV2UaiMb4wKQIULhrt4jxIYHmAToylUiKOMrTOc/wibQZ6kYA0b4iXr0X0H2xyo
rYdkqEbfJ3HrRxXE+lQZNc/xmiyo0FB3IX1kHDIaMkzL+7TS+BPd46bKuevAAWIndkOdWjzTzB5u
AmBRyQ9AwaGRtNap34/ivHM3KYsNMXnGl6QthiQN9whjfZMt9HG60iJjV5p8ZB3zuJEXtgQ+lSU8
aaj9TNAZwR7jmgXkZkwDWqGXejlEiPT11CCCPspcvlw7nGPE9bzfDjLRBFZNKXFVLI60MoZe7aTc
a+9YNylWQKHiJLHIrb584X20VopNsdgLGASuS2o8wEqPF0v629UhyIBm2gLTQ7bispEYdUjVx7C5
IatP+9vCZpulKY6ytAd0j1tpNNhwcuPYCOL8inQNYIpCB1hhCUjuTG7tNTsStUjqbcFnwo7Sxwo9
Umck86kBOpt+13B/BfW8LtAbpJ1Yz+iqTbNWs6UnWWc+eINoxg9JOOad/9U6QPX5ugcOJBxTSU+l
E2AhIpE8xTp3CRYKVR6Afb1wy8Sqam4TioiPoPVpqfB4djk9b1ctu4uwZ+eyQt2DVNf+dLxukLnw
FofDB3wqNg4nuk3GtSxGfwjDCzZ/6N2bHR3sMdJL1ykAT2HBqEddQKwkY8laeYeno5ggcL2C8isG
Qz1NAUzLkEMXKUs+ImGD3wWjFw7fWCigqhpzSZR3DY7H7BPFfun9VVMonRoAVNcf9VdwCjrZLyTh
NmLL5KCyH05S0Jc7ZSEU9Juz7vsaffv9EeRn2fRKhu4SZwlKdWgwwgq5S+G9qUnMIEf/gzPhEU33
yGY8gYgxAjn+iSjZ8cECF2RmwgeYbyhc6xJx9IPhGfvEqNgPjsfe8BDGp7UvgJrz21zVRuossajK
uWVe9eTclaoU1WHKVxC1vbS2v8l9vcAAhsmsxQ4CtE/HClEyYjSGXAS8Tnjni/zJKdT49dYc/+WP
3r8bZbA4e71IyAJcco07lMS+MQ/1lyQxxNFgHGGk7bF+KGWIaNjl44HZmentWMoU99M63D+FAlRG
Nnge+VBtq60JFVzaLl5V9AQyBF0zBtxZk4olK3rNvBBtCGXBZanGtdRCkHnJADjAEFoV8lB7uWhA
fDJWc6P7ObHe1EwyiKNowGT/rEtUghGGeiiQkyIJ8AUlt2qb+g8UdqGT5/4TGfaDUX3XwObdRnVT
5aOzfFjigFRzU72XESEsTvj09BpY2BR0H74b+LjahgsducpBuoG8OgjOss6T2lAlOvBT51MmdcIh
38c9EFcLiqUT0Hb4G/MkdlpC/ZWRY5Z9Kr8MksmvWGj4X4rFX+DHJMNHz7aLvP7bp/8Mf0zhJ0ab
hBf3/fIwmEbzZY3Z4qbrg30Bf91+4e2Eg3iroqvaKY/ETyXPUSTdFWrK5YeOZ1pDHGiluLXEI3bw
ddcZJyH/Rf5UPuN6eiS8fLWDCOt1+Zs37xNVhFm4Y/ziKeeBVv2gqx7AWi6UabwYY/h6qWngcjAC
/icleWsfvIZCaiSuGYjSi7XQ81uMrwevDLj15QLu+ktsPBVV24aOlgWxl+jPA57JeDoQDiFJSK4R
7lqTvAJ8SuenRjpeXmETX98+me3bW79Z067W33A71qOXC0YV8Hy23QrFw+2IVUXJT6VJGrrW8KbL
bdwV2LTPFW0faM8Z/TIz6DaD56rxOqAHKdxFBjE4+E6+oZGXpRU0sJWnrwp/wlEx1XeGxSfBZxFr
QjFH+XDBW+ji+FQGATxkG5JmeU4eD1yrXJ0FymP3ZLpT+Zv7r84709xGWuE/wYQ377gaMLgXcItP
N4pHDFcJnCpcjXoMjMFQB/8kuPhiEmGdCHEy5XCpy42qgs7p6WJHmnkNFXBx3S5SWbFE+jmJ0cUd
OKLOv7xFVAJ/+8CNYeVqX5Yw7sIX9fYb0usBwoRfdG4PppvAZ5Qct7+YxAW1IcDp2vFPqvEAlh4O
Xy+NNRPo+ZlWzfrfSg1vSzCdNf9WePilzJb0PFxY51sa/lZVcoeK9vOLLVdERIdhpnn1q1A6kOrj
qPM4U1zfFnuTr0zS+KNqxrQfgBE7dUeYzlVlSsMgOPXcBOT+Z8OYi1kSg64y/h2g9qvOmgkLLS7g
L2+6AxSNPXJ+LX7oqHbGqvUBdjMVEvSiShyzY9U8w4vBPmIKpGqO68S9Te/FXhqffJQi+UsJk+e0
lqt4clQ9eWWjelFXXTCEOoKjEdY1o3kJ5cGhwYoN9IM2qawlvCQmAcnncJp45nt1IiiWAYMhkPD4
74Jq4yN44fj2niap53wx3jYpYtH85AB5XiPaarNBqwvPEDsHTma2vYYs0XhQoYYpqFfiufkbNruo
V0N1yU6peIh0/YZXlKz+NnZRboHyFZTuJNpxdG1XRws6PrX2EisernRSENbF0j4yQ4xVXme6SF0Q
42yOHdt9qiogXFSIrnTNTwfKa9DeQitjXBrTjVMl8qpWtE38TmSzjby/doZ7XqubNgG52DGxl+0B
dNKRSTMHq7Vbcaja8YIOcNoEVpcVp0hIBfUHuO8Vim1U376GKDPhrPdRf/q6hqh3kQnBD40rlqIs
3iEALadJ6BLgv+4LOsN1MCe/xXnG+jpSQWjHMG6+UswWFJj2MU+qnbg2YVJ/ldUEg1IhsvqJuvKr
SpgxI8upZnCDTlZLkNs62Sqf7zrkiDpXUdqCXZyS3sdckl5h/neMgMx1D1PX5kq8rIC1U3W3QRdV
Hh2MhljcJxz1g4+vPxyn8o8sS1ryT576g6Gg/CNqDv4QeQuuRYpz+gF5paNjQ0lu4mbIXiALh6vb
wzUez6iwvFfBQdNIXUg3Nh7c36SUbhALWCbklkWtWhFCeMCNF4XUp3WvfwZ9M40xfIPuySLTxAuu
UVMxW+ofKBUBfRr51jLbaXMUS+mrvdWFemKVzzkSkTrMi6UfQosUzIKLaYN3viDIBuapmveCNhUg
vETkQ3Gf1VvqVugJdoG4VX36FRb4CrzOmlxSJdTeYxJ9r8QhUdZvSxAPk+V7ddkdA+kXgq5V913W
s1zMpoRPQIgFTVd89xNa1XRwAY10fJqC9FS/0u2jos5dkwsvG0jMVzgB7jkDBm/jckBHxegeZ9uR
52o5LbliovM69irf/yrkigjRCrl3AKyfuM+YQLOjJWnX2HPL697MDOAl/kvN5gXb0D7ISJMWm9pI
U1s0tmXcWWpNKdbgRWlaSSGK/DMKrGC3/I0C0hpUJQFKadsz0FYGU8YqYfWVDQQueqNasoEa/idn
lW56ZyLyUal5Z2YN6wiUblpcLjuVTDq9ZFUYzE/EqNpqG2ua8Q87E0E9JoEO/VL4hqWbilGkBmAP
+XJo+hdXkkq6VTSXg5kVNnnMvt+f41qnKRul53YDBk4Iz8zl47Yreuuoyo2IRVCK0VP8BDeEHUwA
URsoWyW5fI/P4HnGwKj3cnvTiSat3lk2rNcRYwzLTanwVo3ppJNTJesq2IEwBCLjERKrvbLWIPHV
UrSWGp5ymdWhijU68yg6YsHJhOxlV+W6BNcn84G0s9gbppOa4z/H3Y7GeCMCDofuH2ySAnc5dttD
SU/vnl5JT79QWsqPiGivbTfJvStrC8Azh+vO2RnEUTF9+acY1wwr9cKoDKfvxV9mJesZ7B+p2lg8
VHV+zB4/k/rPzolm2M6h+JJk73frtlXVqtrJwaja8zG6aPISARzSsF+3RY6uQMWAg4B1DiEoWNxN
HNMQI2zwBgT2XsmwO1ryV8uz6UBpIcITSio/8731ylHnyfCknFcpNtw+9DPe6yiy5fvMAYnpFQ3+
BdAiTOHqrltPJsteCFaJxyHml7RXfALDNQK6LRFeALQBRYUQf3oI/LBb4z56I+9TC2RX60/+w5C6
w9+6+B27PQq0sJFBxLmA/i068FNpEa9bQYdkr+25xBZnFFnY7FzmDJ2Jmoe34H/XMf2y9lC+uI4x
ZBWm0oOUlG6cw4DcK9I2BADhbUfVNM0LC+KDVWV5SLzeifvXhGAgGFQm66ykVrR1C37OzpvsqxFk
Z6NkuVVBMCR/v9J5djppqUhRE/T4QlJr2GxHjFMnLkDsPPAWs+g05EsMWKwQkrqxQAMv6nKXETYp
41x6+BOGLs8Fbkro7NwlTA14hxxGPhG4fJisU07JzrHmug6lZNHjMSmpPVEwmv0h1cqBkH7t9OAd
MVCaEOv4UFhFAKuWFCxasDlDpUQmneBwUjcagUmRLNzkoCcG8DkLYpm2Mz5CnXoNZar7cQA5MUpY
IxBEvu4MAxJoq0GzuveWGZdjw/A8iVspRHzLQq2JrLSX47fV2UE03XUJ0h2W/tTVxZFQm4GEc+wY
4TzaSgrpCxZrL/pvHzYi+jOjmgjkXn6a2yPjgYoajSy9oO3FwwKERFdalCJC+Ud0tOeoIxeJythj
klqtH0TknWg7HuJrxLtROTxClQEC/s+XR6yqN1KQsY5hBA8fYPjMIkdtAg8JSA8CIWk+jceN28Zf
1Ys8ak36qaclE9XFJhQh5qeyBXJvXSPgxlwMtQg2oMoqXOBcgnXEH3rwjvTL7q1Z0wJclc0HqQOd
P+eX/crcz5QLq4uRepFlu+p4N3hMAfC8+rL19Yl5I+WlXbQbYJ9hwxjrLJQCrKo2Ev4SKHfv2hAI
QVI7g8c5djq2lyfAbeGYEMQAN5otSWARRySH3AYZMceTBjnKS26S5FXSmyEWKV+uq8bHY95ux0np
sFwJ5aiM36JFckvx3IdZiLGViDNlNQ31aoHSBF+mvlNxXn6+OMpKBhgRQBf1Z3FTdpJNyASZz9yY
hzDCoZ5ZCheDthV5Dxu58fmDYtZggesBtg+woVJGdP2e9CX4+VEg9Ormp+W3VxYpTCcSNhb/ihyr
gS9zs2L0VbFLXc9kkgaIoqgnhOBikvgtiD4tSKuPa+TpMsyO30Lxgv8uJuMEuZT/9tbj/cd10GvL
I7KW53mZje9KJemtbMjD4AwxlFwuyGtsmHWuhv9ePmxDEAhQgtFRNez3pT6GpyOzuKSKfOc0qzUb
KnumtknV5rJDTrT196CMK7M8iZGOlcVXQpKdJm7+YSYTWsj2ByGR6YoIC0Imml7vQadRyJPEjaIE
QwHyuW9DuDnmo97QHikNzmBPslZpQmR0rhllxKl71dNTHXvrW9kBsve+4IkUFdJ3rzbRjdF8tWL7
EFyXKbE1GhiG+fdWSLsmp5BoHRWQ5F8IgcHX3mZm1CE8BOZ0QQjMAsjpMYG3SibsvmVvP7IabTtn
ii+V2ZFbNHKebZKmtWLvSqDLRKlLnS9O5o7mXodd2x7W8yThMwYyfHosUCI+VvzZcZ0M7Xp9pKfN
ESsa/kSqqneRRk5RKhJV5FrLd3TzkTuzIsUhEKtKqyE7HWFqm1AOnavzJmHQyg8vgk+7y+iR3apb
vpCyWIRyS9RaHKa2THpo4rShuf4LZcT1Cm86er63N2v0IqXsME2RL6kytFxcTMoaSMoCO+MuE2z8
TC2TwgZUVTw+2ZB1KlGD+L6FKIB6tK26Y/D+8sOYBRYYtnQs9llAJCGPhQH21EF/gDwQRuFlXdeO
pdimW1mxzR7WkJQeeEaZgbJp4YM7B/kmWdTr/wGEH0Fh0XSsOxZirsAiyOE/DzikZgrPTUDS5Lxc
NvrSBiM2RItjL7Jtw7zz4q873ljHNB5Xb8GwA9xBTLUJ4avCjyrpOQsCYd8ZO79If7tm+jeFjhqI
SWD33rlRIJlrWDe4WtOs0h8U2YUZxuOcouYOZYbk9GW6ns3Qw3Xg0KsCRd9FmcUnAAMoE5UYsY40
34N2tWG8dUbreuFZscQ+PUW8Hc48/U6XxksxQC20QkNsTFJFQyZw+zhIh0fmCBtGgKnqZJC5CllU
SKfe5BovlUicv4yaP1eGtKXfw3zictvA9vImlOebl65AMGIZwHgxJKrTaAa6EbTo75tDnRTuhplq
I1GVFVWNbwKdyRvUTAvWh1P2QBwwIW9VABj+4tsuwhYw+q3JtRz91kjC/oBCQoQ500yLH/ipg9JG
TRza4uNbBeWhhIjtWPj8bbGg6dqHFPFKgVE5IZjRHmiszoDbgmn2Z9W04AneYBEOCffuVtuOgQF1
rnhhw+hp7eJMrJr8szEmVsYU4Eaa7FNWWd3e1VWFIGbuVLlfFyd7IXIo0fsjrVgEXU3EChH1oC4f
HkQ+7mTYDsUp6XQ7rN4EHSMEIcDFZ5R/yB7CGHH0A6178is6LSYtYcxyu8VQEKNKN6RSTwZmfxsw
MsN0p7qwtmKrU63vu0B4z0oeRXyQoZEjddvn9ZHidKVVgeNvcuGD5/V9SDOZJ1zYjO7LthYYUXg6
MSxrUt3i4YX4/qjhAu7wtneG0KJTpkxT7kBB8hx/Qu+VMKCz6zjLGx2WcKqAOt5vdDvoVQ72zBet
Lw+4qwxwfXX5pWqWAIIyqHx0XykTu/33iCEsnXBBoZggBqK+i8qIcxVwlACo/7dK+3M8EBfY8DKB
U79io+XDzdOgqOcJaJk+VPrzKDT04IaClv+9sZ4k6CpZUriNYi1YhsT1pC7N+uMEcPz82Qn/34fy
ZIJwEkjQXSOow0hvOtxn4n7Lv8ZZJF/HGhPaCLe8ChSq8XwGjBEYeRruwIQr3H5zGAsHPd5yEu7F
d4Gcvy3zVNNlEFU4IXq80gJGNR9QWXpDV3BMHExJbWppfDKvoikBZOg+ix33JmBiE6gjSS5uKiTx
8nEM15Use2x8IR3Q4ygXCXOiF0DK6Bu78EsV3szMTExzVe6H9/4bid0qnZU7SaY8ifggByWDxhnv
eJGe9cjcPHF9zt8YCe4BadilpITysE29CkYQqHo1Xr9Sfs+smzC93OetSZPh0Z4QCKE3rAovA/1p
fTtRVI56n6V6cufcLGi2OV5ssTD2cUNdUfd4WYXhKEZj5JPENpEuA77c4rmAo2Jhi13f20sndaY0
XBph+GGZRvOqEPr0NmJA3S7E4bbTCjydJJKCUMLuWH00XEoaFw2rbsYZ6IscU/tTZshU3WefTQEJ
5ZJJIldfjFmXQTFn9YMBzstekjRrtiPx7ZWUY1VpLRKmhpWGtsOiumnByQ420akJETIJJjL2hKfP
wFT8923J41ep2v+Dljj4nDPQKJrBM3udMsViRfZjt+aETXxalTC9UrpyU5dzR9z21qfW3Z6sgvBj
ynnqwePTDlJHSkDOsjPiftLLTktowh9T9jswWBVozLZtWi1v71zigrPQ1mPMS+EhYKoIrhj4sz0F
0TAjdWnPOD7DG6/egsfv+peJCBBgc1KMYBYcGuHMx6Vr4Fprlo44rYOREqM484dQbUlaopdOf1xU
Vgz3G5xGIBwMCQ3sJYGD5x32JkQ0qRUr0BCJIWD1ToLX0OLbrsV9/V5Q17iGethVAElelGf2HHaT
9sQcxrQJUGFWVXGqTKZ6Hfy0xfp7L2fUpXkjBVWpal4LwO7u4wW+6iy72/oWjU/YkKpjOOld7ZtN
h1VYQouq75Nx7Xdr3ysgeUwWyAUFSt7tm8XXZHhNtWI90LbbTDdHQDBYQCm/LANSJZQ4z/tvs51G
Y5YIYwkttqL9Axpl0hndcTwH4t3KmFlTsnLWzVxXA4/4kkSB9Ajp1egT5NrLpwPNduyRW1ZYdW2K
kMk5ukB6WswplyfVA9gLYzt917Bj2jI+kjXpOoxqF6C/SLfRbfdggSCZamYgQh3L7Ly16f5IKuTo
rCK5NyAZ3oJ1m/S3smPxf3OP+C60jg5vcLnEWc1dZbX0JOLJSg9O7sl4RJR/CRvTJFQrPzWkdgjf
79mg9WtBOmBMPsu9yblF8CKELWTCVMZElNCPBGNX0QbEAwVyqFCc9xI/r8O9GWqpIwRTx8yaXEGk
KkWXH+tEQIL/vECQRl481NSKqdFon5jXFLawDxmhNH23u5lsrStmcbcGOA9PX9mx2QC2RcIUuc2F
0DzJJviBAznwgG+2t1JCzN8jADoR4lcAWaB7tZG/8MCbJoRiVPpSMPyqKHgwJtFGXa0RLJc8Xhx8
Vu9D4zGXVkbpfJKcP4PhZ/oEygS3WxiiS5iWXQuXm2BT1veyKeOFXGgNwegIGOEBUJ5tubWUEFfc
SDOhqPvH5IxZFW4G4m20pijOHvtbjtECerrYDVImcJahFe4zwctdGRomVo1O6K1WjSnqSfzjs6tL
qV+yonJNu0gYCsZXD3YOOwf81h2avS0whqiV5Iyn5cslUCjk56l1tEmRHC7Fw2IsRYH5WxCUjR2i
C5JRH/DI7K1wJv5Uovb3RrsUM8rybrfJOim5tun30jsMilO/Es04SS95Gj09ccmBF7CBJ/o3Ybgc
Vmu4frGlrAVHuYB6p6kYMfTZpXZ6xvgZt5ZBtc7aTesN1sQmXZy/lB783PUWpZd6ZOj6htTd48Zw
Q7e1wMDMUbOJskLMLIPHSpeqskVEn51oOh6wzaPiYNz+smnZ17CnGtcDTamw6uJriJrsThc+Yw8z
9A2GMtYfBLXDjIcoU+FkSno1ZLQnOAPzdy+BgyhEhE+Qd2eMqvXp1jr7PmpZqCpJusRzAkUgKted
x1yETJlAl9EeG6nGW5kwcmcqOM4H5d1a3zc73xEvM8BN3Hd19rfcJWqPmOnf0Z6zmQzzD96uluKJ
fSXwtZbiUSwqgNdNYhPwIHBdD8jV6GHRpWc62/eqDNdqSyygW3XZhALkzdhCivAGg10FHxdXYf6s
76FmSmF+ghvYHrDjoIisJgIKHYIVfBNiysfwtGmN50lMEUzfAf9pD6CSnqk3T64e4Q52cBcDHbNx
Dp/DvlwzgAvWJG8KOLncN66vlZ4d4VuuCkA4SHLctKKtdLFmaW/AbcXEZgXKk+yNmryS5PY1xtSB
JW+lngolO+KYKMKj/jJ+JRANvh3ukYa8iBR4s8Iiui8v31E+zWyFuWdcdI891wHbfEjN6av1+Vis
wK/zp6qXzUw7xtp48Im7YJud9fXVP9RmZH7OT465jd9wVEy7W85wdZkTPxmi3Ly/j0uwmnis3iJw
yg1wndxwbEcVWDcsweSY5C0Elrqcki10V+FWUMVxpyN/83NCWuARhqkA+jE4sAO/VkUZGJVrAE7F
Uj9xhC5q+VqXZGoVTf41KdE+ZCv3F48UouP+9SMsYB0M9vDMfQWZNuUuU2GiSqqduuFI5QZUKxe6
r6cLZt0MdXh7L+6AWsJY/eY8OB03eVk+Ro/ni3Qdf2f5Oirm0qiPAqd39IYRPHwM6xust5AT8JpE
WycaD04EEoHYTivmEywizrT885JwYxSzaq9R+krvWK06+gjTNaNmhVDy2g20tMTtA+uhPTMNg23R
iNKjmo/vIno/yZT9Pf/kpKxKWUfDhp80y6onJZLwUDzaIjAcDnzqTuZUYXHa0I0mgFicQ1bJdw8v
VpKNSjbeiFPBavbgZw7wJCqajHjClFXQBiKTLhK7+IIJfjjfFf9QZhCmjrKESmdHfXQ1IOgTBLto
1M6OvBx1zzw4N79jE6MyV547bKk4aACfG+KJDPXQT0rDfgykJVxHBzqHEVR4h4jz1d4Uz6UExFBf
7hwwsNQ4rkxaNi3noBFcBdl3ThjKmoP21pvSampE0cZkCePNNpHPYvyDt+C/GjGWstyCGp8z64nE
iaB1Vrbh6YQlXwpurPEvDAgnR0jm3OB323OTHqksiXr2xXNlF5yYRq6KN3ayIybWmXcpWctZbTKX
uL28gD1uYltDwMNeQpRvadFVuH+JHQFnd8jInSh3wYlpqOMBvhQdQo4N6BYdgsILNhH6VWWhBGv0
DCtGvl0WfKYln6u1hlOT4ArwMhWYk1bW+eWiDZdAInLv3MTO4Jr61BxEkncpS6mKCl5mphx9ejjH
MjyV0oydLfIGveVhG2FfbKCAkDdewxZZpdC18PXPOiBdvLdjcdmCZuZpsUC2vkoppBGfeMjAYIQq
hhpmbekq9nZXvVTuLWUzFjMoPCr3ZRMgbLsnK0v+3r8YicBIozqFCZfQSKMXNNznGFsEGDIq1mqh
ZcGsKxKqV1Zth2ehTXqYwKAfUTkr60kt1e0VnXylwLx/0dtHnn+WwXm2rdEHtrAOIDZK7M6ivnFS
/o84AbqXPV19gqSwWMfeoIoI6gxXUIDDnYvED6YMdwhMSxi54LGKWJQc1pylASQPVD9nngRiuxB+
p0FqWQHd3cL4oGCyeROe2vOtK9/Kbq4Pl3w/oZdombZaTyfrlrqNc3x3J8xrsAnqJzRCj6ZVsgCk
lDVHBb1d2VUoNGgDOAginDhyha5V/eKOCsuNx/zTLhUrdpc/jMpFLByEVozPqCygT4I5unWtsHTo
VXb+X9HNc4TYQswvUQEaZgYchjvqGapi7NgYngtOKoZdu1X0d+zHA1clssk2ru11DR0dfYuXnSJT
nTIfEoIgHjK/I2g8uwlaCJdp93o/mF8tsWMI6k7vZjeU48U48yjPtR/vAoQ8yBl1p4ywEjdkTe6n
0p2tWoCYzD9VMQ5vTa46sx6Gzx8qU1SEICbNQ23VFXjibp8tQxKdA0A2UbtSb2p6mf2hQnrXHQwN
dvEDvn+LmG9gsVEW+pefNctaonGBQvKYn6njbg5Hamgah21gI/vVPhUXlzORugsWOXwqprcvaZ7S
Dg7K4WI82zoHC7XuDwRCIKLzdSuGUI3fH5SVyTKm45P6w/vJZF3jC090t9KzYJM0NranhbfV53Sc
Gv/O4TEyzwcqBEdRydt0Y9+hGkqfeHobKCjdinkCsm4q8I/K5vWNWbN6EGtAgw8eiXjFJp4dL0o1
BWqkmdB/nPvHdvD7XDrZBS+dlrrd5emuoAjf4fF0u1AcCS/l76npH9T/98OseLfX2iIOFvLH2NFR
edLRThmT3NYAFXb9PfSdrP7pseR77tQcLGpvMCtZasL292asqB93Q6zdjKVCEh22khvHZAnd8JHa
qj7lu9NqdKMDKauSsJnq5XVF9YpMdOIAKNVmwRsLU5qgIeB850KzaHOSNkR164Ae4RC11WpQMUDU
h7rc47aBXEueoVpkUT56lp7q7sb56VMku/blYGADQUtpct8outerJE4Ovxo7hfXWFxTp9ywqdidv
oZ6CaS8xCfFvNk6D8xIrv8wSbU3MeRyrKOnIlC9F5l1YnWPLT2lkAjWwZkbvdxA/2UATCODPielk
5dwbUAZCRWWMsbkGO/nYFPs6cs45CShYrgamgQ/nZCAFmwbjUjzcU/kYeMAOGs6ViSXgmHJtLWRz
qxRIxKu3H4QVFGhIp6BXBUEZNGIKVQif2RltYQ9EsyIsQu8QFwG6pJmmycak/BYiE58ugEFPqGUI
5OU78N1Z5MK8twRUi2CKZ/Cds3yr9ZXPYvZocB4RTqvCQNWyLNElI87EBoNgmGW651zg5UpYIxdt
skx29IHcRLFZi8cMUEe5F7wN0Sar3lQU/FBYyQiOtkrIBPG93UNiBkUBdz3w1bLwXVtLQVY5K/xS
+DqB8g8ju7+1v8dhnrWPv7RF2IbS7y8epqTR/O3v9Rd9thqcDrzZZNTeNa3og8MQMsudHddKB6TD
Euocu61ozZh/UvWzVDPuzDiy9dFhddryPjIV8HV7mambSdJC1yDtwVCRxyEHRdGkyHaIthnXoFka
EUx6FanjgiZ4H0Si+1uoNMCVOrR/wRz08A5NQwbNINobtROlkNlLTMKlw1A6Lxly9Cxc3SHf9HpY
9zgiyrDy7epE0N+4fXeiy3iIOr/k88Gy6c21+CY560NHD+ApdgJtX4xxa9Hu78E0bD7JP15gxlPG
S3IAM3ijfmeSmTXdJA044Rdub28sLC2U5qcsVWUonwjYXEmLXZNWelXHbtRro/H/dteYJSgssRp1
az/g2RqE6gEYpPoYmCR4ISG8q/3yzPMXookHlD++6LfXFcORcV36P+LTZK4oJZaITOSrQWtInfXN
UA4MEWo58nLefZOqfJnuvvS5meOmOQI//VgwoSSfYuYUuND0uyZ4/S4P8/2FmvY2OMpdK7A+H1CJ
0NlgzpbMZw8hubpTT/f8WT64R/WzK0rYVLsr7xPq6e6s5X3DyAjiUF+fnEzVuZF/giuZSFHmW8os
HPaHYcyacIBkzq2va2Nma1KL9SFfQYJy9z5F4VBok/4/7ol41accrpYp4bvdAd5IywaTqJvS5FBK
wetDaL5pqpWTegLpQPnBehM8nycYbTTow0resX2YiiG2swHTgSGsYcPo5uZ9G6fLoQkYNcUJ+2F8
pbQUKsfD55QorsomC00cty82Ml0KJXnLWg4x4Bbv21aCS/11BUp7SgxD7jgh0XYBUfYUvaKe4xma
ouWv+7nkVsyfe3GxPV4nU+GnjQUUlEoCsNSuk4AZGmiDTbaFKOR2gc9wcSRdZwVp8CL9qVtZCK0M
xWD3QssnGiYs/xElluCOqZ2xZaaQd+kAtexCIsuakWQaqVTMURfkIhEbq3vRoacFlm1BQSbq97Tb
y1QjV8JPsgEDwv5Uo/estLo0l/i0jhwoXoFRweVNAmtaszgA1ksdqFrxgrleRuFpK4o4Cv17Dcv7
ONRy4lgZdyxz8YYBeYfs0KL4gyQ9hd78QRLpbZU49tynYT5A/hMiAo0WuWgIEYppDM0fD2dH/67+
pwboMzJ/szTk/Ep4sTvO+EuyzCidicPjuLE01VBhO4vVjq7seAKwWbJpOpirAEAwOKaGfQVvJwoL
pJ7T+lU68dxCCztRRlC7qWUOeorJR4fmCLylDCIsB7j80GLZuTvl1E++YRsd+ltoxxxMViEXT76U
txKnnFEVvjSqGH8gQNmlDP7Zme+m3dgcuvxMDkvbhR3+4f89G4zAiAqUvownJfzm6ISqcpHRsKAa
t2RQPwJboZldlv+XleeOcN//COX4B69/Ny9oPPw7vKruouBWf5cfddUKyzU7CX+A+MD+lRLaShYc
i8eREjqlc1dk7bJKRDeIIxN+Kxf7LfW5h8qnad6xpK75iZ3AIE24+3K4Nh8/v+mhNvLSPmkdlFZR
aZdBfmyuv3N0ULcW4BSYnL1G+z9KkIlJ/bgK6SrwTPKkMJZxeBvWiKOigMCzlkNq5j/MYo5E7S4t
f294fkdu8xQTC0Tezu6G4V3xk0B6VoymHd+CG0avQGMJKwKTzY6v1xNcC1vcdZaJBAhB/AjW+IcC
JeJyLY5gnKlQIJm+5Vsb9B56CmxfJ+s3Pq4XOA9Uj5re4sc15neflfdfkFngJmCwLzVEM8qFmdxy
0CunDMBSatw6MFnDFZDCYx44RsS8WcXi2a5XhAAQ6aMjX2jzQBopIfNLPHCNQ4/MZmqAmuWTqXyo
imGKYP1HmKSa6kNlYwT/oQNYb8EGtiCwUeH0L1UetXd/fO6xrOFxS2Met0XYG0/kBGQ2TVV06s1a
e7wGvlXYxVdnTnlpun0oVLtfFxyYfpVhsjBn9Ib2fHbPD0+yVx53k38E+Mp/kxhkAiPbXT39Wwxl
ILWC1C2qkCj2J9jykX+3zgi/3hVC2QfIFOl2wAC/2H3FOmLXImHU8fOrmg1YDr6a+PZ+pxQafELX
qwFWYqbOpPKC2iTk6zfSSMlD9Slvs4z/0sRFDp21lCVJ/KSMMfI35Pp0pgANzCS/ERgF2Gef0IoQ
KPYvjyNMlBKVHm3MXJo4lVHqlzwNoNaKw7oyZk0G/U2UeF0vHG2Zumw3mwnMiPtnH1LESv7GhTaT
mD5KrJ9O3JjuDJ9xPz3yeZB5CpEc93TPXobm8Zy2KPD2MfEh2SUThbErCck8GBoMIAAx+jjEAdlk
uQ+yoH1SLvMn76nPu3ueEj6qXMDoFgPBR0fjorhUGhEJqhi7r08D+SpJi79dn6aIqyJcz2CbEBo5
QZpD9ajTqkUiP+lgq2m71LLmc0+werAwl7l77WzXLkJtDLjmVFndx+xKEp4PBt9zFNiMcm5TlyLt
ngN0oACU7T38nXqAJXKivY4ipqRdWhmg82I3c9NpFw2Nwpxu/B4ulhIfz4zZhkEBVhyV7+EvqYYU
Nr2raEFCa+SqgOtjCNlgQhLdeP3sfO0+bOPWqTcYk2+nEBupQairTAHsST1h2QyF4xjEnm1UZpkp
iWyIag6dzOLufTrR5ByLop34Np+GMSmTTYs7hO8og2SlkqaepXRLqG18JQRhIEPQtWobLGxIEaFi
7veGQX7bzzTJlcHroE+tkCO7a1bMvXQkqVGmjr3PPyg3GDMpKwKmCw9h2QT2AQHmCO5zVvsf+vm9
hBO9SmBA3kKVe2wglxC/LUj/zXZIF6b2GroFsziBGWV/gp8//FQjcCgcw+B0Qzr2JfoQUgN0gpZf
SmxTAgnir7/iQx7CjVKWkoEow3gun7bMwvNM79Rh6z5CZ2oZZgiGUNYkcAGUSgr+g+a/BrtD++lI
8RCA4PIWJ9DydrTLuLPN17AnWq4ja55fPK6YsfdMox2Uxg5imneARUasVZNci3mS5N7I4/tt/k9N
mD+n5cHNQ+lPkkrL58LCQ4rw6BbpO2/l7dc1cNemqp/moNwjJUSEBgIZ1H0h8lE8Vj65XNc/1/Rv
4f6Q3sAXgpVnltt5JS3BvCIGklqFLKq88BXFFG28UpL2272r4MPm+hYVxAYyvg0X9/7k3sm31Tf4
0JybgSZKkDc4O+Dq5UDaHvDzFEpIKtrBK1y2sYEYWVQBXZj6T0X4lpy9OB9qCb5gAlBCFYyRT0hH
tqp5WMB/xyDJ/4yauf7IbHo+2lwvfHnpVjmqR73K1ENf4TZZutpFAB0PCO6g8J1TX5xg+8Un1GA0
z0e0X8RyGTseo4KCD/xawOWPj0xkO+esUERJVnQP4MPGedChnZ3bUfW7F/z6bz0pCvkj8OXhYcfu
cJYEV7iuP35n2FM6kGC7NXBCGM9OUiAFoUT67gcCUbDOwr/6YZMVs90Za1bwkgJI/BN1FJ6LokrR
FGP2kJlNQg1UII5FoPMUjnTQlxQ+V3eSyTAuCOMEVVz5YAsrKIsxKx0h6F95CzBE2gq4qGN9SglD
FqAzOXdBclc8L0kkL5C+hnyP5/p6Cc2KSQX2iBKDpE/DVBgbh8nl61N3D5kRiuL0QA69PC2pHAJZ
Up4Y/K1lznAlIoq0xf0rHtdoM6UZ9Bt04IDkCYUafJqDJLjMnxY+IE8rneff7///GePTAivPXvyK
8X7qbalLKAjOWLsViA6E0hB0n+tdXq2vkmBaXBgUpoR/YFP4GiIlYJZdydPEAXZ9hhMQ+lVhZM8y
Yv85q62OXnYnKLwf84LJfmIBeNf6B+KHyuCyoElqss9DPf8/EvLtLJQe3g1+Zux/QbHOz9PkLamb
zxGHurLEsOjvUagnThoKtK8f767A20TclY/ThSG0DIJZJfoBMs+EFsySZHxcwCktoKqhDyZyAU4T
rIZnWNINSP5G89k69RcCNNxtDDV2BexwTDKIyw9HJqUv4aZ/A5FSq09rV8z1WXiV6+vFayQloBb6
xwSFCjk/3/HJ5gAlvFwDgOnY4vn87wSMPsi1RDp3GFiL9KdWFz2sWC6Q6s6W4YQG8eiZrmlubK7p
JzLhOMBPCQhkUlASkU3qWeZ2LZ8bHyOxdDdvqlW9oHBmUkz4TAlVsf09jILtv2dkytnfDIAsbb76
fuPJA4U37WW24erEWWNRer/ENz/oyKU+VkMNhLE6yCuvxpC7a7HuTRgoCNiDxE0is0OstRgyqkaA
SHcF+wX+dmwbZxTK8Y38dYTyhZXUJpyRIBJunozPS0yP+aec56elBaLbg3K18cwAGdooDcsle4Y5
tV5NmQ+YwSx8Vwe25C2C8YuoipFGg1AWMNpyxIPX2GcQGwJn1u5buZUVLtoK/nu7FSCAjBnJX/WM
vCqVk6ZjD8xUfbmFWlH2Uru5ficXRHpkHpcpmAkv7rX/yzEWhHBnV4aYf+3jQH95kMc2HVdINIg8
emeygSug5AL+633HDJQ2aYCT+CQ76zeaEWL0fWNszB76JKNXsOcUdhRu0K0yDwYgfK1ryQ91jq5A
6WBHRXPNY8pb8IeLhWO6Ph0ArbkcbGojPBVYfVm6m0SvcSlzO3hNlNi/bHve1icxOrGvp3jPz9sO
juB/G3eR42+I+jYJaDllSDn3xwFSv0bBd45UGdbRFSrRzUd4778r+/F/36hp5fIDK2M4oquR7bDH
J2xF1vsOAgQiNPwcxANfzl+xlzyP5aWuxj8Pdb9Sidwc5kUj/1TGK9QPmogYDoJ/9Z0kQSev3iZN
Vy+adkAdWjW+wH4rgCHH7HS92HaTtoDaxRo21Or36ulM2oVFqJdtHKkpZVRjNXIRc0LgPacy+lFi
srr6Ir0v8FTRWQbmmGvWA5GT/QxDG1YL1QNyTIualgcgAkmw9wWb/ydj30Wq54uvmhRZxH8qIjli
8niEuZ4sP6ZvjWeLsA/uN2bqnnrp6m7X89zpqY6vZc6Ml6M1QH6EkEmPlkr7hLkw+zvhV5PjiMZu
DGs3pJSPzEWbC+X5a3Uv1KcBshK/1B67+MO/LIzrASi7TkHNbRlXwA8xjkXZ7Pyyyo02j8AAwc6P
Rid3B/Z3RH4JtvVuDZEGldAAJgfO2t5f+3uI9Q+CD0QTrJfPwww7jjlEGkC0qWIuJUAbTQ5faU0u
zBtNhbllNSqRIp3N6hPtX5LvErnxF/DBAP3PpjxBMZzMYpbHwjLSFge621h+Zw8pv0Zbk7YwQ8y8
x3Xk7rld1XqfZsaQ8MUVX+rXv1FmqiB548bRgitPUOZclTb3lSYAEwquPR4jnXFp0sLQ784A9GGs
4O+hDmgQuccgi2Ng6wO22gE4jGUGNX8XTfq7ozdyG2sJbD1x5/EVlmocFBP857K1vBcaG7cw5osM
Y3H9I6m6OBbfVD/WgePpwQ6LUU3viLjNqa17xgGh91Ulp4uUYoz6McyDTcMkfssSY+oEXU7xmi40
7PUbsqgHBZ3V0mypSXf473Ov4di+boXV7duoJ+Wdd0q0hwvziDM2jcCuqZ8W3ZxZYrjTxyiG7t9d
sqoTzvNS7+Dz89ybSPCNv6zqUlsNQ9YlhJA1uCN3zdzwWWblaTJWmuu1LOPKI2F0+tClx/0+7cQi
Xltcyu/m4eRjOobv7C/OmosNXf40i70nDyUgJq4bCTr89Xq70juWP05LJYoWiNVFms21jl+x009z
LdVkQdEDvrnOEd+B3NfuN5mqfZW0YOvtiajgjVJF+0HCp4n6Z1gaJkMbQ8B1Xb40Q0weLVUTJK38
t0bXCoeVNBuI/621xAJK1CEijDXmTpCqillFRCT8JHhcMje7Ymgvclpsq5Y3DDz3q0Gy8Oi3M9CQ
Clapk7E3DC3IE+kgqEA+wWj4U02Fpl7vLb22TMiwajR/8vWOLLCdGjnEKBp34rpyVggdHXajHxZh
r8CMngtH1pw/5n7arc7nSI0neOIEXMy9F7RAzr8ee44HjCiBOBlr/ZQg1K4yK9hodN+8ND4wXg2F
3qGPJY050k7x51B5ZMXz0YBfQwLNZn+SgskTd+4G/n/Bf8SeSQDV4cORQB+SfXdNo1QOzogeMlU6
IEULVGrdRaBOTJ2YckBo/pK4xwnfA01cBQZGOnsPSjxOhI8e2l1wyVdJlykAT1945hP1oJl/ouuK
G7zhek50ULmq7/AltPChM/y0EHYirgy/JBVBeBW80rCtcZGC3o60pnIemW3BPepfJKhWUbp9kAJw
UMcqavApm7wNRe5bstihdPrEOnb1MZ/LXGfNIFhsGeM8XPtjS/UJiANIp5GQav+Qbl/ogSLIF4xx
avJl8MCxRDr4YC8lP78wWq9HbrgZIcUFPIoWzZhlskxc8H3ZfLk8Ql9OBeeJzn5N4QKzO348SBEi
aM9sb9ir8HVHy9FJE1AH6xcQ03dykQR4M8FaFtXLeFHHePnoAlgaEAGDC6DMi5dxOiwPHuMEbIvq
n72mf5TZaL2/EhWdUnx19qdAP4puzXbOker859yM/wXjh6X35It3KiXpsgo/Z14lGKJISF1UTKKh
SW0ElU4ND3SADyPMlOt0ZcxzCHIB3UYeJ/3zMPrfGEPbV7B5TFKPUExUMOEfn1OEw8sNqsLT211B
YymPQVf4XDYZvc6o4D3rE3ifsZrgm5gd3vXLbhfOzjUFfQYvNURr5uaqWqu2w/MizUjhgqA35+xM
qRIgpxHq/yDimlbClg/C7xEQQZFTuSScI3hSws8ZfVK60HJChXPnq74mMdOuIRunuRGBfe8Meq4K
Flz/mKLu+kYOQL0FsSKtUYdBD6ooPzxcezWDklDjfbR9LMGx/P4FfuhkbmctDm9MNQZD+yiBN9o3
jO1eeXE2BRiq0heTCBbAXoWomAICZL5zXVE3+i195o7R7sxnc94qDmbtcS4bZooBRIq7qLKio/Cl
uarcv3omcdhCbUz21Kh7MYgGOtBt8ljnFU/FD9lmyDhYtl8+LzM8WmMCQyhtOv7YTFIK8F7z2LES
X2zzxSTviNuln+mBHijmJPP8pVApbAeUU72vqUGBuQ4oDj+zSoWbaLoxWkfUeQ6EVq7sXwxHE94L
DE/HA0ITO4Agbz65F6SgBORQpPfxyt+kENukIlztoTLn9LnioLP3gppdshq/xgtjhQxITUhdVvug
JgsneOmtie3XdhAiUE0flsXAfBUoOqYRn2noFOr+C2qzbPypNeJvn2xmkpQ292tgx8npI8Ue0p6+
2uKUpuWPeyzkFmjnyfq5W5Dsyi2wX4V9dQ0E2qrtOU0yqFbfU9wNAZKMmDKpdCc0rz5BaCmRN2wq
ueJ0gi0WEzeTCiyT0ggJEwPhQc80FJ65wt/FpOT3eCw3BP5jiGS2WPoAcH2/wzvGORjuESn0nodG
m+3iN8/8qwH3oGyzPFrCcrqi0pKJF1gKwqM+enjRtfO+F4HKX1FCKDLlmFGtNhE3lGhYrK8QIOYb
HrPuK0YVFPn2ZLcl4TzLr+1/IWxZdr019TsJwH+lhy9ZodY9ZZpHlVaSHPl4c5owHvScEzj3UMw9
9lPnyQ+7PoLipWsyEEQaiLJIEtAuNFRZTXoSMQyAxQ0sMQYCeec/CLrNdf6B379nDj32wQ8YHvZi
Xvn3ybIPmvhH6Y3hUVBku9PnSro+NOn1+3U7vSsoUenrIH5RpyAeiAIURW/w68lrUY5ffn7ekv5F
HEJpeJuBRmydx43/rWW9Jp2btViik1bGZ1kT4wQWyt0Cmxdz2VqKqGLLZTJxcvIeIYru0ZQlBkEE
K/VfeDGMVJqIb93lJK+LGyg0KdPwMhFiK1kdS2D+gQ6+aYrs6QyPgIsQHMJlY4M+P5D7Z2oRw2d/
9m540EOumtCWyRlaLfvLrtEvpdFEZU4+9ZuiNIL8zu74Bo/9/G6ZmyHZTaGdkRifpB0EucX+x1RM
akunbC3zISoxxAsJu4hjQBTjW8Snn3cWlU/XT1ciH5bM/IAkaiK/EpMjTfhBcED88EHtdUwFrl8n
P/C7nNInvrDG/d01B4ALUpLWxtyDmYv7/bKfAdYpM4auqFbcyoJ1kL3jv1vAM0aqicCaX6ERZaUU
m/iirSq/TvD0g3mXB5QG4VMk/H04MW9K/ThZV7NTIZYKXCqApYhGeKrDaQgrzKf12frn81XNU73X
CqpjQmA58fijDAY17gLrsREfxrw77Q3Uq+Ru//wmzDhyOYh0ToSGF7cJfPUe4Vh1PLUk6UCBUf6Z
bV9WvrpZam5CaBr79XPveXdL7dNjA4ggj0bZ2J0Nekay5O4q2jILuBl8cdPWVMf9lgJzwBfCEWDi
RspTjtL9WUo45JI+PkOeJ1wRiPs+wRE+qNBSX8gCt9E2CPCnwIxW1NeWDMx6FApv4NsRa0KPNW+w
sY2E5F1M/Km+ZNlXf2umgNmCsH0EPAHshEYJHnQHsgLrGNZo7hiKI6iAotapPAYUudNN/ovo85vY
NZz7BJ1neVY8JISJLFzz7r4vZAkJgnQ3PGzso0kN0EK90A8cL8ESqeC4GPmX2kz9RPcmzAWGTzDC
KUklbGMPMBXmUDLFpTGgJ6L4AvmzJaZaQdtQaUF1qBv18oY/2vduCsUek4GKr0p1NbcHBAVfaHys
2P1IEj04tUUu9mApgsHM87Je8zdygc+2I79/NCwld5smcRAJtIFOoUkUCj4XzNAf3oZYpgUBDqf9
q5+or8M/1klTkg43N6IGhjM7KWydgBmrwYV8w/9jVXBF2NsCq9eVnFc+SKhSBrDRV5/GbbQlOuiO
1U1glqt7ZikNIKDu2mYatS9sFeiwWPqhBxk6OWSK7al9LJAjiuyhfUwoblYY/YDwF/z2bxlwYyHX
85fvP5TXMjXzMiOrPr0Wg+/XEBFlL8UZSKUT+58gy9iDtUda4m3f6xXlADLx2f/38J+io2XN1vP6
M9OVirtBEiiifXRpI+X5bmJWU8SHzF5Tawfd4Y2gRzUtel2f9VS68QNW9+mqhLunGokNklLDKLLy
/+bAMmwwZPdLPw45gsshX4IMnYvZtZCAFF0rq38sA2xN28/2SgQNzLtYYkEuzsUPhcVl3/tDN+El
uoUP+g1GBkUzxGjQWA8irSjsWzXdKy19SSE6VOnMTkTICiXja1m+e5xt4vjzpP9gyOQHuAqw/xaN
TydnQKUvo66CcTivWb5euHE7uoWbe5gweooY1HY8lK+NHMfkMh1+kOFc+r5ct/hq4IQBMPLBUISZ
Vh8VndVHDdzs1q3kDDQwUKscDMz6QwE+ms4UYIUw3doLc6N1kuNuNR4lO9LaOITVYx8sVX/tMTDC
aLokF4NmHwO8xlut6B+Qmh1sRBEWin+PgDM88IEKkiwC2L/mcBtFaNASUwYA4B6vnv2QT62lxUO0
epgVFpyEu9VCQAxqPThki/hZp8ZTAqmfCi/oycCdZaOXzIZG7IIvq9++GjD57MtKM9D/DjbHYGPg
u/vfxFO3w03S4spcWUH+e7oU3Du6ZnSU+PtqzIPoadinMvwG3a0klAN/x0Hc7xO4w6bVvE8C+6Gm
3nmdBcTBsm1pNMdSV+X2pnlLJo/jzJC36FqGxuJyKoDAKo6ZOKaWlx0/uzBMUvIQQKRaPnBpi6CC
yUsEdR6R61JD8wRcA45iVEBUC7UCYClMhAWe3VhP3yB5c7Y6TSDlP/4hkG+HuP04192xYGJbXAZa
rEr4ZF0Bppy7lZd+QvqI2z7UxAEgO4x5mP3OoA9RtzFQciHeNi5fDV15XGjGHF64OfSum9xY9H+K
hJQy5dg12SUGu+BTIU2sclhqRFAXqDVABifnlxoFh2hZI5YbBkEabz4JeUNatJ5P6qc0FeCI8TVG
n4J0CokXCN/smPGUVf9UIDc4J3MYpsOeL82osuTDbmQFVR7yYEhhwdraX5WI+8v3+em1j8mzgMZE
oUviSVvBgP7VoQ+vLtR9vSEEGO3hPr572fygOC3EgYlim15Mb4Wn5NezIHQiKdcyS5/a/N7fmuLC
dsABBVCFudp1SkEfpRBAZIs0rRgBIbkZlk08NJOxJQ0x7OMZ+1Jq4a8m+oMKhsC5w9vR5oHmkCLa
1pQtJElmvD+CgI1tVA/2aJgyJv24x/wfAEF87OTCJ/rniGGncxRs00btR0iuNW2Pzuv1bbzjdV0G
au2GN3/rQPSDtC4cS27zL3NxQvy6KHRZ3m9D739pfVKnf1jZ2GKrYDeXFe/gwJMp9Jvj1gYNnCV+
5AVbVhdwLqJlfosv3CAkCBWj4eAV7KeDym/DMFwnuXzFR2rYOyftGTcxmzSGaHdLA+r0QLG6uKDC
S9nyA+tm346SyMjC0nL79CyI1pj07BRCKMlQtZRpgmtYXsZlhd4rfvYfPkVVWbezXji8QcUP5sTr
GbHtGFsJkMd+RWWs75SkRi7no/rZlE1f+StE0HpcXokZPQmRlWW5zUy5j9pS+VeqEGo9+MqoNMyw
Sw9BY8OFif+DrfuZASNWEkkLdaGl0DRIwgEOpRps0ii8g6+uzZ8VBu5R1r/k8alIy2TGFMAVIhE2
/MGatD2IEdafe7aBsH1qyKHklB5aX+3YUeG5vjF42eyGJ83uo/7LX+/uKNH7msIA2+wAUKMQ1LyU
74tmcY2EymKJE8Z89TKGaxj16y5CggZJs5lHdPrr3fj5HpAF0YoFTNOImcrZ9hSfxR4Wk5Yn7kiw
S9ER6yazN33om9BQIAAnS5GjlKfoaSF5HPtTw70tqe0BhGcAJ/BEQlGmfoAF6o4Ch8FLk7XcMGlE
/5/ehd1kLRy0kh1y65gsdpU8wA09HroVChAwbhM8hwUwY9RAD7E0cH7mQ33A2BBfcfdJFFIOQy8I
W7YqVeE6iPBM9ZZavTGJHQmmZhpysA4Fm24j0x3zV8IigkScQ1+jOtuNaUYlxDnlhLO1kT9Z+Mfg
bgITFLvkSNOYyuM1RJVnFXXZuhHJ8pYgGZP3IFl7zXiG5NompFXaHaL5uQDgesdGfEBnMcFKpFMm
9RrSHoiNWMIheQdEBHel1AEko/lW7fHPJDT07nBNKcXcPcdNF5rrEDkuxt/MIfMjttZAs2KwoIme
SCqBlN5sYyCTF4v1meVizWmciyVWlsbqjHqvUaeY3fcF0eVXdmzPQaUoUD/qmtBhwCI+5HbCewNY
eah7/Lxg68Z9VFWYL2Tcb5FblFgAeeyXXKy7M/jd+z+rtr0p2NvpUhEudtZOu/GDyEElu/CKrM0h
cjw5RiWfTB474xbxWI5C36TUGat4p6XWNIGYMv0hz8EkgEGImMK9PUiQwzjpon3ThlfzB91qwTJR
JnCn3p8R1stCZ4VgZw3c2e6oBDXMT43vD/zvIjod3NSe1ke0GtPYISF1rRATnx43w/DwfOCCepmI
VVRK0bDi5XmKQeUxh+hJEvut8R3IV51E15tV48Pb1jM7e8WXkEb2hmAYqNoH1fDr5qGN43TPKEBl
gTj1s1UKLzo/u1IfuvDCfnFtZmfoKefh4gSHfPy0u0WhSqVUs8PlsBBJZ9g0Km35aSA87Amn+bev
3jel6JF5i1j3UZXKtM2WmTB4MxtgQFVJz+JXIhMfNGAHpxRj/7BJzn7tbkz3sTK2N4y+n4HAX1If
9NyezazR+ApsA/L23PDZ+Ch/KOtYgxoiEdgW+j+ro545JnUORTnqDLjnHRroo3YBdN3izHVCYRIo
ZFMsgWl1yBlPQoKnSvuEHYBo5w23pvfiswLcUKHu1R0/w3gfh0X1nvOAUsg7WZxRghVVz0lxkyPB
6bGdpCvzx6StLT67P8ozlzP2BWhdoGYYbTVFGgs8doS9O5fRrz5BOMFkACr68prpJ9csM3nxzrnQ
a3041r7AKSEcxvm37M6Sy8s8HSmNxUdEE4LAkwTg9aq3DIvmCr71xyua9DQgrPVi72Y0LDDBd7sr
CKODicbdcY9bKbPB78IbrgEhiSN3xPNOCqvrhnwF+dc9/NLl67ozRwC05rAEPWyOqmlsOneQbei4
W8eJcCzMQ8oV1TiatIwEPWX4zDjVh39jxfcDuOzwSiYzvrBofbv5uFf4MLfKaiyqFf4Mep+2j2CE
UQvOzUgKZqVFN4+VkLeu1PLUgWtyXcAarX8hPIgIczsDmDIFjCnPwNMtIdS+gGL6ydomX48g5/dZ
JSMhSbecCpTyzSjAU8eTUN99MLIb8FVJLbsk048UK+5IcJuabVIHxT9VM3Nbtvj2DdaUB//OhAT+
PKT/ajFTVPj4BEYTHL1IzbIk3+yeBzMVU9xs2uYUimczUF3nxg6A8JTZuycgQPdQ0daQHc6XnakA
yPCc5Da3z2/7Hrx46AJgQc0Q+vzvGLsZC4TS9ZHGDhlF8Pp1pq50OSjjMppfB6YDcACdCay0ZTlk
idZrNRMubQqBmfvJZf4jnTCTmF098gGaqZs7rs5AxqnAy+d5IK+74H9DtoKocEfFL8BnFuo0M1rr
dogg/jsejXV8Tj4Q94N1IB9U34wUuwTAV2VpWSv6IhN+60Udy7Iel4IWpiEftbi9XnGFvs+AH4Ch
mN6ir0hfFy8VpZ69D4IYzUIjiMPFAGA/nXx97YQhfzfYNQh+CpD/EhCLOBRBKKPjtdBtu8qFDJZf
7WF1VN/AQ7DdE7oaBLVFhj+46t63iYcERkm7/dGBoLMKF1ceIO60Ai3WrL0k/OO4UzXsvT/pHfIB
jAOdIlNIAqwB0Yt3Ou0UzEyy3TlQ5uS6XOWnB9JSAU4afoliQH+iM2tm3akD8gtDq++V+zcYvD2p
V4CLdKpg63wDDrd7ACyIUJQl2WcinCSmA+2cfrsBqCG2YjWbhYiWCbKQzsUbg4dXnvDg75eQMfAg
xCvzyhIYwRqg0kG983IocYhltQVKUbvkU0Xcc6wKpH8N5HbvBGQefkisf/NDc6tXm/HIuMz0MxNX
rbWuYEy/v5+urxzGMuQgtBlWhgVmOd9NNzYx564TquVHx7Jsq/BNRrOyNCwYY6/hiM3KXQguSuxr
m0u0JfMTccI2ajZSPtc9HYRsD3nFekqOkYDN1fibCqIRCsdsFLekcD9kP/B4dm1lzCpEoG677fjC
1EjwBEq+rKnAoLF7UMuBN2WeFUw4SthsQO8sZ/kiFqpwNJRB6CaKFW1DA/aueoZIo/pAGlWmEzAO
K6F4eqgsWPWXGzoh5Xt6SaulbEktVsgdhpL4xqM0MwwLQEGlr0Vb1xmm32/qKX2vubw/BxWZXPoS
98EMP/igQEbOoM+TWdyYmdbLYUDCZw6TgymW7lufDFwXOMojTQ2cEs/XnNEy6uRMuw74zhII7+T1
keVyVhywjSyxc0bmG/Zju0Ibmv2yoQj1CoEIkEJZNqJ5XzVrgWqTz2VUZTv6leel006sZADRkGzd
OElKGURA7/zdIzkrDrr5ai2bIFMi2jqmA/jE7NGwBKjr4TnShkJeooT2X6O6kgpR72NBqxNRRcP+
Thug0QllB58rdmYXhkz3gRuFWKspjwCzXGeu8kpg3xsgqkNU73vpRNOrfWZg81OTzbaFNsElUmpE
3zLiwhcYOBV5yD4GRFk5XeHltJbB7s++mSvI9vdXp3/OpTb+auZuvE5zgjwANPGovEXWjPOw9TNw
L2xNYXeIRFS3JoMY+q1zl5LvBrK5xJjDQpX5gKmEykN/vBDFg/UPMGD+zHpxah08J894JX49OoqC
DFuSqL1IoZ3n3rjT3+5XdmUI4Gi4saGQf93grxf1vRsme/1qWLzJa/EokAWotXhBKDS9I4AsMbqy
snL61sdq9EnkUo2sYACsWNRs1aWRNmdLs7cIUYIQcxB2+nDvSLp5BSWilMJ8wCl4bdwAuKT6LBac
D9p4qC4vOJQkKNVCPEa9K6Ug32R0FCz1tKbyxyXYsef8/TLRtvfHv9kCOSTCMI1Aj1Qp48MLgKrr
w9WE8FsJ9d4AW9Z8b+0dKVgpnlR5eKgmi4puQ7Mspx5wT21XWQMVxxTEKxIXMLGyLV9hHFrqvyET
VJLSHro1i8YdR/T7RnEx7Qx9oL3qVTAEXuSjcRTaZd6ziX+5CK3Xe4P8DyO1vPJS8+q+NCwLvC9C
CuL/2p9HBW+Z4ig3nFLqHctwZHkb61+d1CgW747zqYWsu4KTOyhAImMHWv51uMVcHZaIEJFUw+UL
/t6+kSDobT4qsN35TwWuqNBYyz6xBRbHFOIIOcfKfZepONNrcE+yNYnp2ke0tCNiTANgx5JCziba
r35HbOn0k5owi0m9Tu9pKAwFzRe9pqrQ/RkZepZqLdx815LYMW6obUHumtthlFu1v45gdnb2NfnO
Mrob0Qr5v9U5RW6/Z6XSd1YPDv+Ur/ndiEJYB5huvFH/Ib3Q/9UJXx/5HHoIX3exO5/c6Qwf8Pst
W4epGyzhmf8nMOaBN38omkKb9ltKClYkrTL5oYjd88yLEtCEBuZacPz1sCeUosV4Tyx8vlYMxURZ
ouzQy2LgkkCZ2IN4uj2HOPRBGKkUXwXg2lXYGIQkrtXUeVcG5plh8VPb3DpgSdA0WcN4kt/Fnkl5
DtCZVzzwT6T8MPMT69BosYyRrwOIUNmXFbR/XGooDIcyW6wfNv20hRtNVT/5lyguwf9wQv8cZB6g
kLrsm14hzA8I4ewSW3BdbUCno7TdfG8mhj6JFq2EOPNbAZnQiYEwNUfibgfUWgAqL0AjgLqwqZh3
DHvpqa+ROXbEEmIq6IFPS1URERtmX8aT7VZL6AJUcYB2lfuEnjr3hZ4Wc30HiEO04EbJxSOkZ2Zf
YiWhZYwwzMFHdI9pV4xW97VyEbQpuSunEPhVenQhWyocozoP1CZOOsLKSbPn8n3/icbye3aUDuo0
U/29+U7ni8l7pMtP4uVH3dCDlMAL+BsWrBxD+MhqG991EDUaAbj05TvlAFuLlx3RAM7tgDi3HNz5
BTEcMwwDoRjRdyG313/xXqPqANoPGbE8UG2QT6vQ7obKVyQO+OKfqN/xoNrTuO6NXb/XYWvDCc6b
IutqC5d2eNqL7aq7t7hFh3umPvT6Z4ua3V7zmB10ZpGHdCH1+6YxzArj4stiLkDDZmWh+rM6/oC8
gPDVaigc5JWaLXFH9rcAOw6DsKZQSslwHES6UTLHFCLXPgXjiwRrAF2xrk+fUaCxKIaCSIaTZvZc
jX4pvFHXNf90QVOjsb2qIpWSmWGUGpw03n9zZ4Pwb6F1UXFSPxiA4wR71QK1Fct6Tw86uGpOs80F
iTAP0nrq75npCpnZc+SNMm1o8zSNHyL/mOZ09HfDR+XM5dygU9K7eLON5gANPFqm4ERMJ6Ohj9nH
pMBAM/rJJwhIleqWAddD+f5Byi9CzA+uzAUWlk6JM0Mv7+DUHTjy2HoPnRC2Oji/XdGnMT/MCQhx
mjY+HO0+hcmGoAIwXw7JCkGsrVsHndcHk2zNNkXUpFhDPohQ8DPygazV3ZwvhMLllpYLjqS3pjcD
f0aD6RL3slLGXPd51zGsbNN198dAIr3+5fQMXCLzRRhtoAWiRB96Z27Z0x3uTnqzCV6Xdhc0H9ye
INnUR/6S3UojmA+J5zCPJbHalWp8H1v7lNw7QUkf5cKbMtBUqv5bKHrT3IKpTw9FeybA56OqKjlX
UOfzR9uRdB/D+QHNcfdRsaL4BR+ZQJU1RxXUYfUYpWVQ1m5CJhJdTUljlSjAQATn/wLG5rK5QIsZ
AmxZf+R/f86EWiYo6EQFzkLtNbTZT9mDueq3UL+s3qJngLMITF11wggF49Hk8d3wfOjPfyZpuB8I
gyV7CnoePVaSLX28mDMDqq+Uhq2rf7pW9ptIzBXChGjVIAUrTvT44DJhEC/1oKPJAOQZVlk/2CSV
pWg2tCXjvZvsZyywi2PE6VWwX1B0fo8bLIn7ATMipfXDtnCRm/eEAX9BjgyE8wI6Hra/RLlNxEJt
wvS7HDlJn0rHqIFWBWWFKA/lHEUEihhD6833cym1tJEtv8CcnybGYJQdYQhBm1Bf1tm1d4e5t+S+
IXNoTxFg+Z8diG2xrzi3Uu4cRCXhjxwb0tvDPUU9Vytuv1ww6/cPUkZBhBLtgWzoJMdHdLBdIOF/
NKbwT/ieotDQEnK9FGDyZxO8dIlvPuVFUR6PGYwMrNzlVQ5jmaeXmyeAA6CsfqWHhDmV4sdRYbp3
HfNLYJuK6f2k1UVUT0LZF+GqukSrl03HzFcPukQbUHansDgp4isj3S5yAiex4YGgr9d2cy2Le0iT
cmQ64PDCmxQH+VtTEn6qVPxj4KbCZl2HPIGbVSbE0j4nSdV+NVzyRipUaWgWeS2cVg8okNWAbBQZ
5OvshhDhFzudzcZr+EPLojH8U0Y3apqcIJ2VRnX2xHL5QbDVFjZSHlGc4Uu1rvfNA8sQTUW5HMtb
Fl9mCWQKgXcKulWs9Cv3/1XyZec5WBHkjjBej0ycNTZg3yxlmfgmoW1QDEEs3d763JwFdo+a8IRu
nl5kByB2aaE9W/SvH9hgaK62V7fS513Mr6z5PYeSgeuKngWl5qbxUZ1X3VknKweXgcQTokNKV7Lf
W+azkur6Ipg1gg1KxdDmSjptwj/gUKu4uhOLDGgDhRFKa2GRrP0n4E03PKeWEsiafFaMAcWK4qmG
uRpo5mEOcfc2QsXtsKiALzdK7LjzMYzEfuwNZCof5aBFMFPiJHkqvFGY2doKQPKfsukgCbGbmehp
p87S4Yjhp64iGAThbYT2D/d1V2FfwjyobDhDNWw5hFKThtZ0l9F4BauyuxWz8pG0xmFQkdpN6/Oa
TM+vk1BhrSOwnw14S9UQOqp+9gIy8F62Mi3coCZIC3BL4Xxhz+rGTbgCMi1ZeDRXEGC6WPByv3sS
XLBZ/0OojmNTEtIhlt/1BjNC8hIKzOnFLZ6+iRoXquGUyWMByJsyaTxuvOEbDEXdjjO5s2FjeTzs
eAVIKHN8RmOMPa86snvq2JpLslgE3FdLWf5lj03kFNftYR0QAWrLt1MywC9Lp6Qwrk5wXU+3FUaF
anmRvBWA0uSVGQPnLAjThAwC+oMKsdjpP4suOpDRYSMdHMk6c4N9Zsoi17qY8FozPrV/0u1gqZW1
Hk+ojlq9J8GtmuySMdWe5H17iOeqHz4DnBavW9t9jHmpqhiZQbfQ7gzudesd+cJpuUudUXUrbdz8
mKh41tcz8MlUzeDKaczGZTwSCquErR8HJ89XP+e3ugfPyYx3EBWBw8dS1u41jDLM9lcJeBoFHo4T
w//sLK5PXXYcrlG0r/9TAoG6NZsI4d3cBXNu2/ELJXP4JKekUD2yBpFaY9MF0WtN6WC/vPZiuSUb
+vZXp43tXPqAXiqFvvvBNf85ISMC9Fer6DP2hC9zkmgDla3seEO9eKgiBjczWSRXH1161VJjrk1F
iMoXPRtaQuIeOejDWEnQ1RLCayTJ6LkLkpDxf/P23AhthCqa/6Jb9tsw4k6oODRPHb8r9uLB4GaK
IJNMOoTG4FXafbugZw64tQfsIS4hDzFqLtPNKGg1OE1n0RDIvDME1P3P7b0QLSjiZZ7AY7h8Vs+M
3lIJI7joVh518vrYv53d5gx+oHuXqO8Vfv/bZKPBfrSqjspQ3ELFUMr9qYhUYQv6OOXLX5HpqMLL
MJ0Op5Pgbnnwm/pfwkkpCgq+UPrue9n9KvWMgtryzSvvcBwJexQO3KjJjI1eZ5MbKHKGTZo4zOqs
EEfaLiJs5rI0MS+vgYPOL6sSerDn8A3+ANIIn8ohGHateTdG5C5nTsh9WT0J9O/T650dKWQIIRC+
SK9Z5lsG2oxbYsy+6LN/ZlgQEtyI1zTAh8EqFYHdmANyGFaO5B8dp/cXf9uk065Xfnc4KUGjirQt
1HVvkqSEKkdN+fOt5lDmD/YblxfuwO3kHOhPnSavixdB0KLTlwY5WYJtjif46gyd0SB86qn0NqOJ
9t0ZOPxCZ7FdQQnN1g3pUX42vkzI9uSRE8DicL6WWuherh7eek2Yrd3Ceuqbe6n1WyKXzBZP+p9U
oYtcY6kWaItioaX8ToX5sQf+zJjPoDf58B4GGScV4eXPWBsjjQR/kHsXlgbbUlbfngDW1OHvpDm3
5xYWsEjXIGv7ldtodNhWHpYyBJKVRbROVVWGlJZMZuyM5oVg3k6vC5uVjYVzrpp4F0Ih2mzKhzhB
NgX/i2qphpPrDNNOIDyASyM0R02WJKCK/c+Uol4ej/NoFQouDyiL8CrDGbMK0gFahLa3AmzYq7KT
6jm/IrsKf7I/o3JOxS3IA6JrOxXAUsqEyLQVNnHZ7LbMQoD7pQ1zbM9Lr/jN9Y0rMJusoUcAeafH
2+3yCXwVvRlCsJXsFUeoUu57XOFCDTm/aZuWzujsPr3Hm1jLJ+/51AFgA2xL87jU+V3sylWLkA6D
w/MP+JG4A+kPr8+SaEREcjoaYCUKYicIbIXQgehj6MLQEftdLe03Nn9wqNB6cjXZ38EvOVU8GmHk
AmMEo5t+syW1/k3vjV99R6WNj0pPzxM8LhgUKBHzCsUUjI/xwFBhO+coHRfe6WFALidVLWUpX6PR
Tft8ZqnLdgMrDw66qUSDDH66WS8NSnXcFExcwSSJGMCtCXe6rIFliBZgQjD2ZY8/HIagzzQUj7el
yfAgvOCdDv5jwaH9rXazADlOSWdbhzRTnPBZwoVWyEbOa7cduTU+UtLNQpe3bLBXNTwBAfO0K8/k
ReyZ7hUJfXKNpQG71Shp8SdJNZNxCZh2p9iusQfQEYdoXjKj3NDmSUc49Qgy/6CxqT3j2MdtPw1D
FKW+hlPnPLSI7Obmg43X79bzgZS1Q645zdDVDoX/zA60yoOLnDOXUMVOyJERmiAFe6EFrS7zpdNc
B3ghNMpXSmXPozfcakfZzx2JH0Y7vb++s+JrgWEOxjdz6dbLhddpGXv0JefMOkO0gp7TieV7LbE4
jXGyw5qnmDtFZwKWudn2AVPlQaEm+R0rOGXTgLmQcYP7l2Gye9rkDgfLEB7WQI5B4/+XYgEld0mr
mPCDCTCsSXlZjyACOStI1AvWgaUMdZzvW7kCTyCUFUxFLy8MshnD2UJDRvADzIF1PT43zKtjolSj
BNTMCQWZhUrbgrEdag2TFGns+c3EWqxm7vCnZwmW6dRatLfUg/oX1nem0/vMnyXv7hwBrQOwKS/B
/Ofjfcsp3uPrJjnsx+smutlmRksvvH0RuM5tvU7zx1HL1jiJPOOsMGa/z/dY8re/gfyajWeK747x
NbhQSgXCtu3TCcdhISythtFllZQQGFkPC61+Sdc3MJX/INkya05965F/l8zjc/IiwFXoLUi9+bb3
B2Hxi21Wjc8gszuc2PJ/e0FNgNuKInqbez+UfqXr6ULmT0lQL1XHV4ST5YvhE0p7ZKPefp6VS1HW
s8hiDXiWyz7ycG9o/XVoWZKHgh6GWSTKc2d+DtB0s2GIEIbBx3BWb8g9NPUqAbABshLm8pqurWwm
GpmHkDXdai1euQyy+oHO+q6PmZJhbcCUYaC23SPeGAArTeBHmQKfgOR6bJawqx2nlwlheMi6lBsT
WvWoyjkbXPJAfNXyihOJZEgp2vK0947IjFAfI3Swl0o5pjSDefCLLJhsXHhNSSCy/A2MHuGu0dld
7Dml7zdf5+VPaU4M3VtEhLH6wN3LJz3RCeRHNa+aQHyt8scfwANYYbTLpKF3Nvau7sMbkA5jd7Zw
ekn2GVJlOEEdL05N78q6A1LPALDp8dAhkAMggLaNC4C8xUzKlRWgsfTjdTyOBX8eSyIGeosd7J4H
ev3dwW2BM4F6sHSCBaR/Rq7g9czlcshrJaE23Q0ul10XDdenVQ8pHag70L21k9Fj4CbRG6b0J94f
m/QQWARF6s3c1Of0h+bWWySJM+PqmvH/vgCXjWs4XTLd9qRU8+uPNTwCxULMgwWkrye16Qte69NP
1gtnYzOkQrrUrnc7yf1liSHO3q36iORS0rxxzUfglnzg61IZCEBNGRp//d5ScmfxS+D0nmBC7fBK
fCsTUNBlPIo0MIIdSbbhJI0/CSubwwj4gEBKT8Fnrxwp/ikTEi1gAi80EsLSDET5pCI0DWkTBGgZ
Rr78bAmp3qqCZgXvoR5mI9HTiQJmN+q4eWXkYh+0+EiNl3/DO0+vmkagT8Pwq27X/guvgNNMmjpL
1mpJXI7p92nj2aP04x/+7fxBWDo/qjX3YIheNAxn1oZ/ED82VjTVY/MST2rcBxnkvHbW1FRYeGmu
DjAgz4jRHIqRqXJ14GZCgKOIamgqxcHFBU8MCLIaZRZjY4jVISU1Kpt7rgK0QTqbFHQ7TnGcXlq/
6I25uY4HNLq1Glco7afqcmYHnRi6/l0F5988ADdUGKP+RezrtBhTaJYd24CJvbPxRPU2AQv5CraS
EsDCjInaTppR7Zc++TtPVWEvhrFAm1hzMDZ6fc0mRkHd3YdSmc1gjCBqUehEGTKhZ968BNXxA/fs
Xoo/quvJlOHfI/JH0NKVxX/nJr7wu8V47w3v/jc2v0n5X8UpnrHiOI+rqWL0WXh87L+BAwSdo+2M
oEoDSj0dAe3FfA7A5nsB7DZvNc0tN5AwcIJLNsyYP2HEzcVQouOzZOC2z4AldL9CbBGIKy4rh1IV
4iSdRumh7cTxYf67q4/GrvwApoUO+yM01aCnuALJ6zPv1velcagWhuM9k03OTP1LGmLEj40OTh6l
q10JgV3frunPg5dRE6jr7A108R/b/nZcOWlCxJWKuBW92rFZFXSDy4PTVHmyMcYngiZ9UC9apICo
vjX2jY0vR8ZKb+foRlOagHgtjRpqST44P2y/HaLVMlknZm4pThjlGCbApYDUd7rZ2ti39v9MU6m9
8fYYPbt1tX8YRcrPYmGT5FS6u+gxVxXDQn+PMEGuYEn67aqTbgm1QDPDIVz/5lh9tB6APYsHR8cH
env9UzGGgLD4LFhhh11zTj5XyPF02/xQHJdGzSeOI++tOet4fR2x3XFXPlXrT2esfYPgHgaKnkCW
eJmB3vfR9mNhGozurR5hF3BaKdnqbLx+GNM3iVnDUfP73eZY9ZUF+wZC3heOrLCKW33dQuyhUf0A
wLs8NTHmIu/CHsOZGWdLdZzCrpMq7uedfxzQBu9lQwsd2ZgqZhmzUnsjCa9EZmzgDJA1fIshIs0+
NAm4JK1zXp1kfDrK7lvL4df6Q+J1/TaiTwAMchccFL8YpNfWHR8I9MMzdp+Uor2yphLEx6vj5TqW
kOlCl3ChIknt6Hgy79tOpdU5UDMyE41nS8J0NWozvBjAXZ27BkrgQW6R0yswTICoomF/D5U1MOli
w9iL4yzsEU8WtF4XEaSYtFDzjqzBg+t8mKS/ZldIoPKi+g8mS171/aQPoFx86BKw7jhdkbsmwmIx
PaxjOPrEuNTUkO49bqQDeMcEpTuL+a2jT0mDNIMQFQUBinKChy597H+u+rErq2XMhuCr29oXC4RL
0FWtyXbyXtxV41ZfpuGAS/mH6/Ba7SPxONRjShit8pT90//Yjka/obD46w2PiktU4v5hGs7vY69F
xg6ZyzS2++BzCfOujMfxMXjMa++JzFOF0EXgxYnCwdmJ9acoMp1mWqRhvGUevWOUNJ0geG7hmyYs
dS1yz3Fb1NRUdsQCU0mJ5Vg/xFLM2H08h3QevtRuTBqaXKPA45FZYnEb2HsCDjZoKmS0rJEJ5or/
J48SzprwtYAcvdWZn9ythalc5vfTiP799lqm2IJc/ifBJ69xXSYizxjt36AUI0JLFGObIjD7uUp3
1NOD896L/o3T4Ez45rkG+1LQkS1Ponxl63oSHrj0NulkvoG2GEzVJ++SzlEDcA4kRXvqs3f4f9/8
g5/JqaeMwe7CGMWux3OU2uTaWnu8N1hIAq2EfIiOPRRpoz2QQ+Gku12ZBpbXBelGKHAqjd+kDgYf
otornfOGDUTTqWX0T3I0ak9mUGFA3yJYLBt9++84V4M/BMXTu2eQRqxuv8tiAWDl7w7FH5Y1XLhK
6r5b+v2INjOIqFMfEqMjQ5tBjkGyhGZNhgVqH4efg4AtqBgRp8b6N9lkxW2QLjcZ2A/vnF4dO0Wi
MXr4EtC9+d4GUkmxLtuFHbFUVQK/2B+9Ry/cJZehBwf/qKKUIRNOjD7QxE8iRb08YsTYS1wmrpmq
3uqKAGZ6lrDWqXJuUYRz2ABtlz7v6B/zhbBjimTq8sm1QOkT6Efx8tRyFB98FRPgAhPyJnrXYcEu
n505/vfA5lN4k3cImfkaN7gghS3Yhkslr/GXkMepYt2pf9Z7rNbM1aN7lW+M+uvHVBZOPAVSwkJq
G5BOI2bWMXhFXKL2ga+KjbF4bxuidtaK1YIi91fl2+9GlYCrKbfTw8HK4egdx38o9L0ie4HVENQj
f13Wkx6sJfOMjxCtI/HRgrXnZ0yI/virQnBOoWtMh3WrK+rDOeLF2zP8dyiCJvv5gzht0PpN+Oqd
Lkxj+1v4TC7crkWwKViTViCUUKUgi29ZulrMPbtftRMAIoLx1Tx3JxhfrdUyrqG9vV9r0WeH/cWy
1Mqu8Mp+rGUYi98wdR8wLISUnc0DCisCGuSvtXv0Q7rPGT3XJOQMxQ6Ug6paKfnIiJ1hzulylkb9
SZttJN/0zFpsgG8wTC0nJ5cdrLXf0gFKIuk6/god+k+9pM6aC/kYhG4ASKGABfJH9CENDwkw4HMO
hzgkoVl0GJ9pcfo151PgkW/it3UXeUnZX90BPz8uvcfCNz/F3Ln2xosYZPgMA9DKWcRXueYMw33b
Im05Sf2kMYCuLINAjSEm7ohEaWITkiMzOFtLIC9bn7Tr899UDk0bNG0xX8Ryy0U23q7DtsgLnFNZ
lNdyIywZ3aMry21sJV2m1h9hEE7z8A3vbJjfIr46qyGhvFK6tnWSW2y6Dq6XFbNk7FBo69/FA4ps
3tyYv2zL1AK4+BQM4kG0FKxjLdm6Y8236cUM7Vb1RipqlalGwtdQiRtBmo4oNuzLN94ozylmojb9
mh9VduAKnL5kuGIR7Xoh8WpcCHp5zJcSf4FMQngCVpmKdk68Jpjx/GdVySlXvxiHJ8xVy0yJ0aUI
w2kfr4EF/yW4U5qZjf+K2RsjCN16i1v8v/8BEcExb7ELwqFr9oEjH0i7U7ikXmXZG+Pk3/QYnvlL
OzqV+gW181CoBHtlniKMr1j97Zv3IGR7yuP27OlkAEzdKPe2nzgajMxhRvPatyDNuNJxs+1fd6n+
I2bYDETa9IV9XEeeRKmqEIAbc/9n4MamMSKdQnvL6VH8KuDUYFPiKWW4wD01m0nNzZ/74iXxz5oi
sUeuyIPjkFBTMcvpQQD42kuYsKShtM65gMg4Bcc5ig6hpwTERhGsKRgRb8fuPKOu65gPXFIrRg7r
vBznvbGrlGv8QWLBuK9rok3FhxvJ2xmnIk/jEw/JNFXBg2/kSb8L08KgqbaCzw0vF6OF+2g05mVd
fbztW1iqviwSOrGx7tK7GyGYqmFkDmuvFqTgm+UfLlsVyycgM2WIJTuERrI1+Nw5TTTWwdzO/gDA
3hGO4RaKq/vd8cW8DCwezFAooY4S2Y8NECaMSqXFnejhy19opaZHuSMV0fF/qR3RqwZC07KpcRVh
DgjK4QRacwB6DLMcbr/R+5AKC1tEdGEAaKjv6AwZfxWSSUmplXCIDGyybOtshSdsLoEJK6thDHY4
sFRR2wGF23L4WfNv6d4Y7kEel3GcLuvUbEht7AnLKWFLG5yCIP3heyNEKv5kADdAxElR1/zxpBMX
xhEAxbT7MqIUYI/OCgLOrld1hckXQNadXdx4CV5LcvMFdp03d4tTGNaoTSU8CzurETAgA8uKlEWS
vsduOXmKun8G7Z2aLLkKvZn7RYvRZ79sy9jzNY4CESZBKFJchL98gjXl1K6P4iCJUDQJNDhSbayr
ulFwOnK01foHPgCYCuw5i7rzQjdbduP8m780JtiizUw0A+KIMXJ2GjbMNdRaJgJ/7Ku2bfMqLB8I
tCyd+zdZnnbikoUZEye4upeb9JxEWOJuRSuS8cpCp3i+6Uq7r+HUZBUOJJ/JFccUD4Cd7bT1Lpu1
mWDiaZpl45GOWOqYlQ9YL1mctRJmcg0idcsblR90AnqEP+tiFRE4aHguHjBIYklp138thtealfx4
6wLcOSuhpuUNUay0hafxp/hSHIy1A25z3t4gYkZ32qqDWLrMTUatoyqPyvpCfa14YyHnZ1Z5FbIs
ar4UkxhH9gOoJhfFJmIPrUboplNcnhlezZHnoh4wX2uOlf3zlZDU1x3bg8JXfCiERE+O3Maj8eZs
tUd5O6Uy0enS5RHTuaDcyvM18JKp6fzy46sZq72ak2S336HGBI15QPd6cUnD0EEpKZdIdNbfFTxp
krX3xqdQN9ajd5bFg+88cv1N7EQ4RSrEaXtN9o08AwKi/WIH/H2a2B+5qNMHMD+hkwY+9pQwgaxY
tfcXmWXMdmYMSp8ZgATOP5n4o+VF3lZNJ0TKTyvUNap2HTlG2enrGJYswfc+Pyuqai1LuZdcovB6
URgEWZL04/j1W++VCckBGwAWUpXT3UadeGplfVeyDxx+h+4ID9t4bdT+23HAoi9AWNw2hZnqADRh
YdE24ygczoWiLikhQxYKrawungGqNa47VEhMShtp1u7DJFVNklivBLgq+b+wPlmUvWWSQz3kaL/T
/PHb/C59awmn4HWFOEtwAzXPoQyQ7/30ecMKAMKFgLumVTmAyUK0sMz5eu3nfGNqZSnBU72VaNBe
IMeXk1ASYGbv/E6vyEW0qA5bsCiwB8iwwn+s17F3DF+Em08ss+QivQOArVLb3MVRo6TR40HFdut3
FmzeR8X5eo1PmeK1walrGpj4Lz6t6XmwZ1C0TzUS5QCk3V7gLGwqINrAxvSC7EHg0lgoIVgYo0RK
vatNWCBrxhVjFCHZc1LN7bLCRkbo7y5f5XPjUvuUnZiF94b+N4r1DdOL0sgpJgzsEFpHE1sSEylM
QQeHBLYPbvf+s4vKe0hby/u1foXUOuUwnhYcHYBJ+uuhIKEyqOYKaXJ+7ftIBexdtLo/oCsB8eRk
7yFVCbKhmmA+TCH6EEzoK7AJV++9OyH5qi3lOOu/T4DqRiE5FPO7q+2iogES9olTGpn0gamvrwMh
8HioJFrdYm2EEbjYwC2YuKVIdMef/IEM+j/DHWO3tyiwF3/zggff/ICPHwckxvaH0LE7FywLVkSc
D//3u1tZrKZ2sus1Ur+CJmNmxqfGhzeN/54u98xJjmVhgxanbWQiuB7lVwGFbiHLsjOVAaBDggAK
/WPUUkhwPVmtg88yzenoayh/Nc2nfW1Sd6ilTbTueK8N65sg8t7V/ivQaia5vKJ2j6Zd6NSE5BEL
K5ZetloJpN4bzPCpaBFs6KBTUIYEPDoyeLkmfrFT2PMo36Te3JU8m8G51c5MFgWx79/7flF8satq
lY8tyKD+69ZuDLXzEROpyaAUp+TjWVR93bACdIqZvkGPzxGhHUhNGrrwe5rkAqNwzlSkEaZW1woK
xGgPaJQHG8MADBamfA4OD+h0+MHSeO0N74PX8S5TwpCZKMxXIGQKVJaJQHdL9q+p6XEMzFV9AGzj
zjxjI9F6nocTmRJw1/BUBWk4lfJKpbx3AXMnusFYOH21CniYDXGxjIXqDxi2BEDtopfrkZ+Nafk3
fCQwiM5oKkxO0e6NM5mvznzs4q8y+ndAykA+D3W7XSVTPRglFFiJ7YaocN0mveLBZaN7fUKp454R
4hzvJUrWlxD8a+Ly5dZ3OwWwFECOod8FSsNRLVGoIdTIuzswxy0Nu+jA3YoKLrVXmslTdsTnD2FV
+RRh6SeXVBLhrAH7LUd4YNgC3yKRwwZKXdvXxEemeF2z+ZyOkj83Lods/TJSQ4hjqvQ/8Q6ZGUOy
lhHHOo6z9SJZfyUKlioKNBwkB/15hwdcUpyswsLfo60LTkNTY1rrl3dI/iwJO0vC1wePWyO3nol2
ngH7wlNRa7b6/Yo+MnyroeLdoCDOzqIJlt5cpAdfJFYDDX0+UignLuNUSFHePowbScAqD3leYH9R
62bOTge7sn1t8CAsbBST+hl2kp6uIQqfQHun8p0YPtdKNuT4AB+qIAXcFtm+l7ZCzaPbtGNvXhs/
JaU1UQIG+9ppX8LBT9Uv9C/WR4IoJXxDBtIk2NKfNZoiHJfVlvq6dm976SGbVV0//RkYnO7W+BXk
j/SR8us40/2Z7b/ObuI2zfsywaru50Kon1ukPFsGWlBcOMn0BJKF91O0oSqXg+G5zaUqm8Y72dQc
4NVgZfFHjAtyXPAxq5v4ebNcOAkoUpFrKzU8iXj/Nh0wI+mf6hJoIHLO1qPkQTvTbxbB2ZKjy+Yj
rVFtM3i3XLuEdE3qMh4x4AsYwjhU6b5h2xWDKJfmLzyJ1x1VCJPjKnEqWpDmZRE8NVKDO00MLHXA
U4VV1Igpxys/uXlNuGdvbmbPsLlDOwJlnkc9eA+Q6GFawg9NNDTiYIRtlS+zOKJv4kRorNRqFaes
8ejiydRSeZUq5OxhkUk7P0NkY1zu0+ImW1TBhr8cyFNibIrFsCtiT0J7/kwKvtXzkX7zF6lzhznB
rHc+BovHJ184tvcOKKpN9yolvFQ7iLZbnfNtNAkdALO7F0WG+q4We8bV4jRz5d72DUM/VEjYwzHa
sg50RubXlb8TOB8u1YxvakU9hnZljuL1Oxn2IRtklX+Vh4nrnZt0VzvYcDB180r1pdr7lRJJzlEI
dQ+Z45j9keUJyo0vLthDLbgli3p+h29fPqf4l6RfJk5Qem0itOeIupei0FMMTmK0VTWy1BB/AJPE
q1fuVet4rcgWxngX0RVxoi08fhcmMpQncdyfEq9UaW34OEobGMYV3TdPxs2tuTfnACL5dYl100MW
RShFzgQ501oVXIdIzoQzhJqYgCq94719JYY1rKYdqjfKsIMt2YNA+mm/ZuGUv7tM99G+FAsUBvtj
H2m65ASSoPwXFTNIwdDeucbGor3/2FtQ4MXFNK/DFYzHI0/uxCHhYpIJjO42vOJMbgJgNM37LrkA
BYZRh9lFyGWGnrjU5J8mQDH7QuOQzBvUTwsOEp+WCnUnMuetWBmxpxBduSao1AA5b1gqwoEPlEHx
3gBrfaMkB97YZJn6YXzW2OSkz1eUoHwmDZBXm8hTi7lLniBQvmMuDeQd6sodtWFN55ZrLpmq1e1e
OjOFWv7Uz/9mki6PxttUbbsnPRzfL99S9gE2Wx6PRIfIBpWTWE2+VYFgPtrpJML6YL0UixVTajB2
ehIwDvyG69zgH5BhnYnCqVbSjCZGx/RMoyHLjixk4UShYmE7PH7rlvQCeibMCphXIRoFmpvuFI1Q
0tNDn5U2gfsI9TWAieIictpxUghs9lqzTYDVNacLvOBDUvxJZDMXca9XAzZmqPKQU/QpkEEPbWrN
Mh69/9C3DFaMTZmP+VZZQGSRV4oqoYuOb4q5JyMj/hw4KdST3LwfIFGV/bSHiMg7DjewJL6+oqYp
mrmAGaP4EDfbR3J9CxD0JP1wkWKTgnyhfPPdbV5crlnfv2ezw8BAUA3VRfNHhcGUZqZFQFXbPPnZ
UfMztHZcx4TLczKrrfcA+aGJMg8gg8ej2DfNYqfJNjCuoh2/yYwB5dle6tnHfCKrZdj2u8UJHJvh
LTYP1f+b9s6Btn/Wmv7mFKC0LWhV6mzd27GIovBMKRwixOIDhRWU/QFI/5uhscTWel5Oro0JElKz
jmH2XvobZMwuFh54VCmOZ1GQztGYGkwVn3v14mcMwzvJkXuKzKnKwVXryhCi0NzBBSaKjFiJIOBz
3tVUQzrxcjXJuxt7i6Q1Piu1+3XlGgIvTT+SFexKC/L/24mR4urlgtK9pDNNYrBKCNRxPWTcVxdL
zRE/sTVuNL7KU0FbC1xPQaal9InKWDqV3aMUYwcPZ9XrBYUNB6jAeivoDSx5Ipdqa7nTFtqVN1V+
5qYTQX/banaSqOCA9acejOgcQN0fAZesUkrdaTkNZAvNLBvbQN4rh6Dugvnxp0IAt9SFWFh7AKml
hx4dgCokJiVbtxXMy0qRz5crb8UmQP5tTCkIqMC3ns3FbgLl1Ny5EZIPhqZgNhL+ub1/rXowUbGc
nUAU0nBqXBkgpvyPR0AWPs+OkIJokUFNcTLB2OUvVKLjzPLQh5a8tGA8TaxVI0XiScDWIhoJeBRP
W8BqRvk/Zn+70Jeep05ptZ3cHvb/i7yzrB02VTf1GkJmH7hU/bt6mE6hNuEiEfqUHdWc2imu0DRr
xWpJvcXVwbaUetYsaKDFarW4GXBJOa+ltvkRsRx1aP5ELYr/E74EWn7M8H9PDpTNOTWyLHgEAkxy
lcLVLb+I34oFp5sQU6W7XpTZnKGA+g3jvdxzE7EDl+j1K8RGD1mV1yGBboG5DT7i8drydpXOh9hd
VPJAKudAJsCj3RSveQ9n7v8F5dop2OF83EkVfThxQT7nkPIZD4E55boooHrKq3W32nIKMf8bcz67
G+YNjGI69/6FPlZPEbWZgKr5YzosleepkD+ck4c+MOWMH/UIN0XC7pO00Bxek6/L+uUSRy4wT3eI
HWW98WAABAgwiJQHNOeDRC1/xHxLGQ6WauxsuxguaDxM0MXK7Yb/Ri8I21Xr0obb/6RB8y8G/xXF
o82gPAuJqNIn+PDJBWkkW6OCxsWV6FhPKU7APXIZQ4UnUHQ6X/mXSb1PDXU+7kO9R8/s5GyQwvQu
3+s6Zdb9+b46MrKfHmzeBW0U2nAVtDH1TeOiKP77gtOVTdqEZop3lWL9HN3S97IQr0papU/f+/Cb
Wk167TO3ikKpn9Yzg1IBwd8uisw/MwKcvqXOx4uU1QNtUm2LaGQE/vLpSCD6ZaY6RHnXqkDUlZDu
ow7YU4HUr5Gyf68S9cDg9EbGKZhTW6TwKd2j8NkFifMU5nF9BWTtHjWXT6+y8hRXEZuyx04LZQlh
3N9P66wADNMB+uajMTNtERDnH/YNLuULNMzVv5nZhfwZJ4Et8pndFbA6YhyVimEEZ/6kPljb9f6Z
raifcF9vvghrXoO6+XUlSjfrKM87d1o+JeCBS70nSORqK0FNGcYAkNnXFtnrRVRALUmMBOeb3Dd/
5Cp8o9h6UprZiSHO6lCDB9qDvGMAynpUDV0AIxR+GKak9LxF+WPKMxwGiHbN/Xuf29MHsnvC/h3b
Mx03UXoB/4hAvwXZ2HfBqPyyOfJQDYFpXbKL249XzpV0dVmLZ+2jgtxVgPQqwHhuavGT+j5/apIG
BMBqkHZzbPoBJyMAwacX2QOys+zrnYgcXZDF8a3f1H6+9TL9TBNb4B2OKLYnALjTBsFDzyYMNIWH
yvEVRbw5lDjlx1rUaYSekrMzn9rwavarBE/Ayt+V5wBpqxGWCnJC1TKj0BB0fHhyWPDWtuzIbMWF
GMZMLhfkpUxUt1X76grBRCXwOjbPlPMSS938Yw4ooReDzEyDomxQIH0zZ5Ywd5gxw9g1D0a2AHQA
7Qc7VzZkVCn3aI/tptr+V/0tXC+IKaGcbPx6TAoGjUhdJaJOnaozoXjp9Y/AANqqu/JZQVVJBtQv
lIeT+3jjphZVySZYseUmNUGt9sBkGgg8aSgjx/84612qAox6HJfzNtMAqKxG+m/1qmP/YC85CPWp
x0ybWzWw5v7mRM/2PRUChYdgtW3autDDO3oZfcUjNTS9cRliLeldj1jGO333S4+Rr5AxC1sa8sHe
DGdeDzgWWIg9RrmMyNS4Kuwvq8MVmkEmbYrWN9P+vp85IK0w74waO7yBR+/g1ggvpyHsCHNLIwTs
A8+XOD5wdiNFhvo7g7QatVoP5jlG6i5czNUXhS4Z/++BJKYKXBxxz+C+o6sqJZKD4Uh7Gzxe+vmZ
8+7zRA6hn2Qgkv8ylgbAEj2ZE2i0MCCawIPvbI1ncwTfTeycyLu15XFZjz+BjYyb6M6stQXKAD+4
G8buQEGvzNlBZPgGCKue1KXkA6j3LKV6lLX1T2C+xhTWsd2RaCfDmd3cjImdr4ES9xa3gdMfyhew
nGgftN5G4NP9uyFMvr8zGTh8JIU7eu2chn/9psOLodepDhCTQJzD9lPBBNY+kNsnlhMq6j/juJ7Q
wVqhOdkjStDLbtv4L5+P2jbFpOg/4FVjI7AcdBlobbA0Wk8RtU2RPtDkP+Kk4ubZHXebHaV6aqxw
fB4ptzgmb7v2cA8jJkVYbneAot25oPOQ4NpBTNLOEkTaT46lHw6wIhrBGIzlzM4DNyw8GWvwY3OD
mu/UdXyNKhxfpX8Lrazo7Skmy0H9fMNhw5FzbtTeOYkeit9F2BrTcIUcJX3bNCn7D7q5/7WPjsJR
Q497TNWyr+XHfx7QYcKDMt815zZvowwrKM+eFjGwbuUMhN7mMr2jj8bCwXx1Hxbr6asXySzRxTR+
bv85ll0TLpezO7bcxLaetKkhy4HL0vrIf1ZSOHEwNfjiEK5PmB2dpuNO7xYOf1CTEw2EC+vTbBzn
5tr/Pu0nKQlFkVX84t2YCsR5Ooh0kaEtvOOFHbBLYTHEp6qKXoJdCLszrcQOr/PW0yZ/Qqbk1m35
LttngKXGxZBJzCXARIztn8NwUXl+XjtjAF0+OO7QIvmTr3lcdN5CBfjrCWZdwtanryqIS77BKbq4
j0o7988ByKiilQYmKkmiuZcnzPXzPVjZqTPPmcKMdVuxUa4Od+NG1v8xl59Y4qQg1dqT7PBcNLD0
bsGivQp+eJFgyPLglHVhC5zYQ5uPKMPitaqflt/QRcyTVAAPBRcs8Tnspjcfpu7s7Qdog9dePRPT
zkSj9GtoqloLbIY++ur6SJrVg4Lt6Pza+Cp2JAeG4tEcuqAZGWIaXkDLrGZtv7f53d0kv933f/LD
AtF5k8DbxsZyX33BbCvoDVzMm1klz1ipCgaPSk7dAs107qhBxjuBhQlnJwihopoLLpiEmh6aknoI
JKBEa7aYTaPo4J24NBuaYv73dEIsw1CxXh2gqJvRN6ANMcge8ClRUCdesTfRhPVD8TTI6cbs1AU1
jM7FuEJ0TSaNkrx37bPiAoCmd+FuEqz2EXFYMM+LmTq3xhvONV6lx30J0JSgnjeV3g+E8BXE8HED
I9tSmcPoR3oLWBbJQke0KUbm68iU+pLu57Oxs9uz8aLhrPnSJg8m5NywSvVhH7ZjEcD6CXk6kms2
LrzMb9LSesOstRYcVKRAkM010ng9jg7TH8nTmxL9v2KAq1ctuZ5/TrBqttDaviClhCK+Lez2uI+A
7CDtWxzt6kKAwTDbYn+vkWqVNd2aJWJWBIaNX9NntrX6T1cepqjc4k/vM4yd6pIodf090HEQbBAd
j9mVkQpfYt8RXAadaAJJCKrvI+JgoXgWQoD7VW2/NMjNfM20sCGKV0J07UMzHZNvn+f3PPk3G+93
ygwk+U5pDQbg4pE1QDkpMBYN6PV+oxbY+0hgEuoJ3EmQazBeAumKRTDXI4N5u02WrpTjjf1JW47p
NngBL/Udk2PeXQof6UfTx6WmU8npdVYMGQM/vpCqMuF53DDkUWWumeHXdG9bP4v6zEknbqNKu5gx
kaFJekX0XGcuAIVQ8jwLV1v2ukiRnxQdYbSVGtBoSChKnQDPCn6HLeT+dQuKPd363d9SmQEjP6XA
Z2nttZPlOttE1sbeHvWeSTDem4b/sub9DkFSbvQCSdLhjPzOCQbPDEISsO0IdQwZEb0y8lxLyi4V
nEx2A2AhwpUfROxGJuw5YcoKX5VXIdxObi2ObJNTbxszK/TLPA/qEqj9ikbKsg/oOxDhwT63IB17
C76ZDd86I2Tzu+tE6Rzh+DwNxQy10dJBDEpaT/PNkfHZI2ecf7PgSzbkuPqQPZAhr+2JbZx9tk/s
e/1fgCsQTZuqPjlVVjke1WvPpUIYD0xB7oFx8X5Ux22Kam7ECKbIac5goHsbAZn+2YaWSkdU6TSX
BvLnM+XZQOBhzyhSBHUhGJ2tkF/zZmovsDjeD54B+pgucJSIkEf5s3AwdJfhS6xrhQLmBS750n7E
pS1DlL+L1bkDn5jPtTqrkwRLSGLnIAv/+tmGaDt/kGHjUVYo4GXV8G2uJ626m2VFrGjFyWm85c4c
UYvmmTbyu4JySsVovC//rYOArzgFRhdNVS89qM30e4cAiwj7/HmzLD5eldXpPbdEkza0mjq30d+P
JnMTZ1+Zp20J4164BJG1lJmcd4PIpOBv6BZoYbPOK0iNAFR0AMUirwJ9TsY9xytOxmd9TTtYDjV8
4nmEuhb2307PVRxQxDA+ZVlBgJMk5+i5Ps/pzXkoL/XKNXwzoKLwhxNu8TTNaZZrFGvfKQPw81sG
MXcwSMN1cvtj846b8x7Rsi2bB2AIbRHhfJWKxEchx3mmSIotuEvRmLFCvVseSca+QjgVkq6pyV4g
RnjJPWLkoph8dXKKc0/fSmsuIxc5hkXENLJYy7XkaZo7jFeAHJgJZfhmQfd48Clntk4p4bvVpaUt
iH7EEnVBCxG6Og6w39NfJXCE3+3taQ3c014SvWF/0d3rQquDoJ97/jMW0dCHPE3qAGuqhvwM3IWf
p8JIbjcZUYI/iR1cdsUSt8iPq5r4Wu3iUNBfB9PWOCnQwlfGG4BxCTPrNTrtIeUfhr+yMEcyv+5x
lq16uhbQIy7QGB5ihFCiUvpaewlSCWFCh1W3y1SrY2x+Au3EFds0gkvqxNQzIV5XjvSPjShQCKkF
Lw+zi6wveotICFZF/tgg6pww6Eaq+8xqZQlgFu4xwPXE4kOYJOF2MkB/CmmvCL2qUZjiG5Yw9Yq6
2dGYqB+WvdaXDA6y+37bn1AN1sFS/QbHfm5SChX9wz37RRzyo+O60eVr7NRr3I28zwsgRKylLYDm
g/+25wU25HZLHmSdCmxzjFhdtIqRM13B49eQTN5xAIR4/sgrRcNICA6KYn4dTnjnkjJhKd+NFh+R
x6w2B/CZ/Yph5+KfEjs056FGRNwBE1eQ4Kn0ZvYs5elzwlauyeArXQ9KT5U0dHqy3ZkFaotD3llJ
TaBrDuFrq88fVXeZ/H4gc3L0wIRgmwHEPpcYzDbcqJ8OwCOW2Rv73IuKSBzgOoSd1NEUDROoWK/5
u7Of6bCKRBx/cn6h5I4XPji0B1H8tZvffQSZiMpPxvKgtHDkgRyD/J8Uj3dgI4AJPRxsSz8A85Je
FsBGIZRzggKW2KVRTFpzk50XRhg2iVBVMa9TBWqLCah2bbMW7M8IM1gaZV4NaABkAgW8kD9fxjcw
t06fjr1fscikv7hzRNV2DkYrYwcyyUCG3xQG5027WBw46Kwn/dmPq27aPr/ivSnJI5gEjG5CZ05i
R5m4CxuRgTZsjFf+KGx53PLTP/B4THrl+tNALuOaFInOV5TYY6AMKTiZT1f4wkqU4cq0PIH/dBnh
kheTdiwX2DT6kF9bWMoQS94A+rt2CVGn4FnqrF8maWT+vn1Zt9RjmIbxfQlmmsq4+7bGyw01TNew
1eiC1QXa209iLf12M3NOOT2R34Wv0IzEFPMNzvQlFfA9MXG25ubHxyiUGFg1pYeJKghZmscLSyqg
Y7tNa+5b6bcRd9IZUj9+cD1zUC0j89cFdoGzxAD+73mTWlOUWoNMYBheEUwFU9l4JwkQ3tXzkLu6
0V4nKnqKdJDDGt86KCNZhJ2ClKjomsD5Jhd1T7B8Rnce9JMPTabRg8aMUgYMlr30c06ROjO7jVAI
8bUoPnFNjJ/ptqHE/BJ9KKWM46IH8Bjax7bgI9bFJRXHTOHhNLWD1onuhNqa2Wu7+U0kUKwaJVDE
BH0sADfjeKJUDVPxx3fomjLr1p/2BPu3+rfT8Gmm4KsYW9ed+HUJhnrpTx3dzLM9/SH/jMEuQ1kC
1ektj9x8J2ntsTnRQLOj5Qlf0LULh5K67mbaZvGwifRJuQYdnvUXIoUDLw/MgmbEG1fp93mDcg+A
zG11KAPc6N9VoidIlYjRWFLx9OUxMd5BTfcKGSHmnLQB4i9pPeNop/jXZHx9Y/NXs/RfAk+S8Jgc
9NoG29xnUcfSuIRwA+lF6Yu129rEBMKCAOtru7VvynEsEar4euqLxa+oiqJoVj+ZrtqY/Amfx3Zl
36WoNneTHARIBwnLXFeEVBJ9575zx2a/sRyyiN+/7/0YsbkJSi3sOzNjTEY6SW0y6yPsJCC+uTQ7
4gp0UodDHp2oSggBk8ouD/Ez2pCVHNoeFBx3ZauOz/D1FgpN37Ncfwx95/wJemV7/D7xs1MVrnth
cEZB+pny4bZZDkjz/MXSX1/R9vK0reiYB/gezoioklzJgVnW/Ji0nMOCVIECmJxy3yWDLi2raj9o
6GofrHyCANgEK9SRAQHG5TZMuT/dyKc/bXGRxRlI6gHnlRj82iasDUeRW7gqbsBZwf8qaWIjIddn
RnDsAZacET9wkXOupoK/R+PnQu/3NkzsV/83854KuIe8maV8+UX+SZUJLXQqUCKepVikiIBSd53R
UUHR2WCDG5sZCrDH2/g5RhVSMhWQ7FhJqjE1pe68ly0DjntbSGjPkTZFixl0KhzHE6b895Hyzxul
CklBb4woJ2kFDDDxNmqLUpgRwDnRI97+QhXy57XcWCnQZqsGo3zelITPH4lAkood8/3ulI9mTaFH
boQra/gUNtBRoxYr5OSWXYq76eQmtPOyNuGwjZO6q7tWs93wWsR+50ZjNgNuNshIuxPKfwK/fCam
QvDPCCSnyYT7G71opxCHj6ejcyVFVGWg7F3/klARRQou1t7kx6qXO0dgj5QvDQUUNxojxm9rbR4z
dx7XNYlDqm+Vu2a9+MH1c9UDMfjad5LWETEpyG4m047yOCeu/0LIU0x2oEeSdKsC6m6L0HM4RxsD
DVjWPNwJ9ioYKGpJWBnyO2AQGJ5VKOV5o4509mjG2caBSArbU2rzK8nEArkr2NmflfqhfZWrWMy4
H+YBBYhXaxediu912Qr6DRo4MpHaEZds6lzL2VvF7ob5Rw760c92yRknrcbXwqCcX5fN0pvgKxeS
gkF04oY6opbJQxxbpSw//E0CjjBUpTpBnGKdE5ed8D3mVB0N4rBWiNVIegNgK/oTC6VS4ghrcgq1
rK9/tFoXBs1158xDpWmdGEVrmnUJX5mHqlyYubG0D0gfUXhCOewMB65JfgNdaMtCAHJuK9iBzWEd
xdb6LgZ4x9W3Q5ZrCShGmpwb+S7Q2KhX0eX7QfcrYW7sNuOsQBdykQtmkipOyC3MhDgxOIu/pEW7
Uf1UJuRSczfrAE0g8rgV/u+MDm/b1szDbleTttlsnjR4N7DkStpD5Tu9HsJuagxeBQ4c1Rbl3h2l
1ddgE9vI3b5MzDFcdBo/u07Pp/iAz7a3YxjX6hetxfWYYKoG+sZMF1IExwQNo7ihmiYu7BfM5nbV
2wttx0yf6UIq5G2uQj/NSr0NbEfAxRHh7PV3fGg2JGg7SCNEbvZMQxy42e88Fa/ORhpx19MymY9I
EjcHN5zxdREJk+KITn5CIlqQSX+7pNsu3fYkejrL0gMyRaBW0CsypUQNncc6NfPeZ+qovPkWp9yo
5xnotVVGmQCOBrISBaav8nO8UdwPlypFM7V3CsDxzg7QkGJLR+UBy0n3GW57RQmPnvV7m5pA6tvd
lnv4PBoM/tI3LcE3L1n8+hCqsmOEH2vfT3hf9QRD8CDtOjyg1Y0hRJzBOO5DV/TjYkx07AwSL5mt
uwC2CQmBAOsW9kqYPog5hiHGTFYRBTiAFUYnM07MOMdbj2A7RVh1YKRYa7Ju7LqEukXQmJIRm3IO
PQUlSvNUMgLhlgm28WohZqBx4+8GOX7FXUbtl9rqiTw4Ka8CYgEsi7wiH3QPMZI2io764n6QSFqH
Ibhsgyq2e1p+wlhCf9N23s1tnE4dBiLdV4bfFh70lXR6S0KshNyrWJQLSbWJ14O49Hwrh+ghUzSV
XHH01LsAKn7sGNl1qla5o104PPeXA7qLl9Oc2wLbgIRdKcFdvez98FIwt0gCoV5yZ3jX3TVdQDmS
rsgZyqybCd0U27de/hoiZgTpnX1h7gKerD1QQprHzkID1ReE/lrwlwmo2ZGCOh6Os2swF+LEoJS7
0gsvhcU54GvFJ1AYN0zrBLp13RP219CA44+KFbh7DLR1+kw2Bn4xAqC63Ccj86vz/BZOVpI80W37
qFKWYyAYWXyDiscRUyN/w2SwQW73NO7ZUGWdFWozILJTvoW521SIluVA84tLzP1F/KF1yhm4K+eC
uV2RbClcubGrIu6kOA5Zoiy3UsJRdDo56pFFqdz2BCFP+EzijifvDpe5XKPCLFty0c8MQ0+102td
jvYNrxm2tHSqH/+sb4nFnwBmqlhAGOlheRgvVRCbHg/mOxQxh20nNwv7d0rYvoqZUv3NkMlgspnt
u0qTbOozAwP8jZlvrOlcU/HS7jXjaIfF5x5QbneA5mqZqwEEe3s7v8dAgJjRjj9uT+Y8hdqcS3aL
OrNStfJTlYbhLx7lxi6JJFRnDohncrZxQdpz1OtHJdxCVc2FpyGezQetv93CpURO+ZvFaRegRDF/
v+IYeINVoJXLtBjvxuZdMt/dL0AvvVtkkeN5U27TUlGQKRklGRHanDeM1pqaCnPW964zsM0eJpPe
q1JXVeJPcUOxdW+k2qKJTcK4EWSUZKqWSgInpONeMllC0Dc5Y37cqvY66AN0Xhy1wgnOUvLQjKcB
npEDmhLIYnfUwme7PQMxkK8IbQgS+pcZQDdOQIoJpVXWdU+l+vDPqN9vajboaoSy9XpZ3j/ww+P8
sKZlinE2mCjopxL7oQbagVXSxhFyzUijtasU3b8++/EExi3WOm+GRQ5exI53t0doqXrlg65D+Cki
J3DhaMzBfIh5qV0Z9QzdRoQmS5+Z1JD3TD3gJlGV+gHJS5iiJzRR8/pTcrNZ+FqEDS8/P2/cCorA
fej6tdrPRYCfVHOTxoqL5NBhV3VezUgjP+pTBtQ3Z0yS7eXg59Bvm7v4nBpHSUl8TEeYej6919+J
609T1OlRV5i9GZHYfNXIrBjuzUjrkdoVdiQyM4PORc2NXhv7pBj5ANxxCSZMuLtA6ZrtaJnAAoTN
hdRcLe1xKfU7jmclfDgLsHfHFlXr1hmMGJClYWEVfTLyE70VdSgx61vGmoH6N69pTqTCPYn9rwoN
t6FjowawvhY2I+P1XmxA9yENniQK9gfXyLj+sRVEzN0JmZYQCzaZ7fQqkYHBem1zT1FU5NQWbq81
1VpYrelbjPNwX+X8Lq+QOOKiNG2YcNAj8T0FyXFef+fdGDi+S/DaUyY1nBDXOPvavin2wb5FQoMU
RTeOYd+8RY/NWefuNKk/p9KHucqpF1fKQG6ZSUO7sqkUdnBHDG5mDSy8TzTQxqEI03zlXNgsWgNX
TGQQdHCVQfpEitQi0xIUMmvwtt9ZsAtzL/SvRaHCe1GPTjapLdZGWS6ui1rBH8Zyn149kqmT571K
xT56TW/+3meoHLAfD7WfJORp8dG2yjKAg0x2jtb7tDTl92vpIKiG76/uRO5HM/I7qnVThnypeIAj
c+QBwM5Ci0S2EG+oCcmonpXX1NifHoj4z/H/A1gSCf8lnsBdY+EB7Ln0u/zglHtaH3mG6c11IXWg
JJodfxhL/FlWzG70Le22zC3F9GpEOSL4ko/WbLtp67ii9Cejoj6HDafM0FHOmTPuT0YrTmJGgDQn
ZSM03Qxr3JyHW87ePu2speviqVXKi1LY0bYq3bl4kpscQSbH6ihJzPgA8fVpEY3/2iBjnWiydqUi
bnmdlAuWkgHXpN/dSKjU9HDDCAsi/g1yeJV4elXxtf23VMYnkmaz8U4TFdTMbn9iQj23Fv/PxPpq
FLt6dvjGZy+M6x/r3YNOd8dnDp6wexWMwkDsqAPBkn5rP4NASysnvc2rkVl7dI6PXXvlbSwZHN3G
t/mjdvgHVsAxbkWoSAlt+lJXlxQhuVCVFAI3loCbtt6TfvzQY5K5Qs2FXzZwNrxVC2mzv8hzgVZc
5gK/ORsYIdz8OQBj0bkhiDArzRc8OkwE2c+vSwMKE6CFu2mSaG2v+XWnrgCzv9irDa+pcs8O39CD
Lbhk5nRyEyZoAR/k3Jrvi0qaG/ODwxh6pMxKUSCdeiOmOveECAph/Y+7rb+3bFM+Qts4N/koMC6t
H/qJCv4SjcTvcxjWicdqdA0xNf8SXkNoI4Q8S4YIU2QvoA7qkuIg7hxzrof4R2dVSlKxvQsdPYGH
jjZ6KldtKgbSUS1tGuaQs0Kwe+cA/rqS56KIvoRfgZGPVHOsGubzw+6sbZSZwaSbAIM6qevgzM7w
whPwjggSmphgB+eESBMFcKyRN2Pr3uZDusX13P65Bsvm0sg6lSkN+ULLZ8+4MBcuMu2wWoWO8o9C
6tElb7mnqS+35wwDhXIYGjolIoVJ9KPW4W4qAJgSjZLG/8hw4wWlj8FEdrrtoPAwegs65pjG03QU
M4GZqDPgUPfcNRIhPfA7ZFTQEHWGu/Z1+hSgmHiCs58m6oVXMoGJkrVZ15zXWcw5jq7XeqUDF/0I
GR4pf77F2O1lHwYYznsbqmbQhD34pfh3zb0vQDY8UkK3LqqW62/29MdHqX9hp9eH9nCtNVUhl6nm
LphpfuRisErDSbyXGRXmfH/V9Q+jG4QYiapOEevGx0vV/TWQhz/liZ53IwT7kGmT5CSpoQqig93G
BbgLgr+EUsvu8E8ipY/bhCo9owQkCkoUowFjoxvDNX2+c67XTaSq+GFbbUtwEkvGCezh45sWX/zB
LDVUxI3FrWRDd5Tm7XTi2Y1C+HZNJuha344rqXAYqLj6cSQGvrcJ1iBcPiNdBuEkZA8pAyWH7FDV
4oH5SorlS3ghlT6yQvB5Ik5azYcTSAVvlOyslc5F1SNuhbVNCOXFUIu5+Ww7xqIVroG/qWszSX3H
QuGwSo4enlkev/YBAMR7ybkME14TKa/m3G1b3/7L73Mx9Q0KYsg4ZJXCaNkdHAW4r5nCQ40hJkcI
2a06goqRQqO2Pte4vdVmizmvxBhGwAsd7Q6NZRewzF3sdJttgDAPFz27cY3RoxcHOrDMHXwiHLtf
r9G8EDs+XZDXJUy+jCHsVxyZHGNEu522/sLU44S2aolpVji5Eu9uy83BjJWVRuNgbpSU9T2q8Jaw
4Qt4XAmClALzAdyO+x+PNjpCEQp21dC3qXDRrqeSo+SHaZI66JBKTzmo92c6KGBDGarxwzqwPrKo
YrD3biCVgKl1hmlyVF3i/0UKKtXyRd02z+YBaa34hMktP2RVScjoiFyGT3QTDTbckNb2JLuuKyPA
f7aDwBNrek2ImFnMaP0F7QwkCwcRi6JNLOK5ADLFzwFNkXd3iYG9AVEDu31n8+cnCtcmHmgDAs1p
zzo5TYKF6/NJxzAuFy8HSU5d86UbFvEjNDzSLxdf0sqGsVTABQrO3Ma3tuO3Wz5muYrthi7AgsIk
8j/Kh8VzTKmWozG8xw2ifT1RqluwKMCXjJQKGlP1Yr7A5dpmF4GNHRBTCbWyap3jeNriRVsDyp9+
oSkgLJsVEKo66aPjnFfqaaNA0Zk1o88ICpTn+0B/Mb3HXjYTdMWDuknXKD7biys7xIRJamUWmVeE
IwvjROhI80hOc7t3x/qwwp+kpPQLvIOZ7gNg2qTDP4UOvLNlRv/TsyOH6lNEzqQFjMvDCwyaaRzR
KZDIfix8Qyqpm9ljZxBmo8N6dx9GIrP26MF9IidxBmwvlx6KH1A5yFRc0kMdFhRkSVhxc7HlfXgo
/KbeYSthIrI8dwRHixCkrIuUONJU0vMtQf4HYSwZ5bAA/+dq52SKMJDkxfUCCxHoYSr25d0pj/0x
+whSVqz0znSKjl3wZklJC/tcErTI5J04ywsqXWAzAg6oXEANdB1fkRegMiLTze5nubvDeJx67NTZ
ReisEcBje7fN8KWFeGUEX1/ceLP+j7KMAQuIj6rACS4Ye4IY6tSV+osQAMCo1o/3PMvQ0e4o62aJ
sPk5EzdXGve9wSMtia3tzufQGbnmSvR30HojCOofLvNizxPAVy6Wak1qedbeZ1c+HKwNdv7AQySP
uzrZdh3fJsayzAm/BOpRIKFWVhS98rmB5z17xNgid1xN5N8QjDQPgZL3KF49QJA7z96p949sXIve
T4WVGi29e2JeuKcr+JaPpbHScpLV/fwByqqb8Iz0jgVI4mBkmn4gWZup9XdE5vlRCU3RlNamHfkx
y+gxkYkE4nWDo69CDRK6Hn3gUfvi8yKNMsf5QIAGKBXDyRrnWHddYSbEFcRvPXLzWyA38DQ5owXB
jTRxYBVrUfqFbz7LdBSGT0acu9aVTCom15yMtv6y50ZAUd8V8w2IBmkeC4FY9cqI04ohXxQWCzer
itWvzoB2oeAGq6LhXs41YZ3jr44S4Z9MgLpWeFNB3cJC8EKToqwjVo8oAIVb89iOhKppcS2ZXiZB
6VQqIZGFOtCIGTY7qZAifWbe46cxMfUoMvmv919YwdW1EsKfHFLonem3PDzl9tOfFvu5ZSJYTZQf
u15Jwd15hLVhllUXSxAnPPwj8+Tkp4ubMOgxot92csN31cqgRdvwmUT0/SR8S95TKOgiCFiDp+sl
tnkryyTvLrnpW7VXP5vrr7AxJOaq4IoiXGis1NoO2RHI5K1b8JNpOUvSH286zmEQkoXf5iNzYhG/
dtNm1rhXJHcmmg1FFFQRcNE89mxMM19Yj/dx2AcHDM6MG6gd6DZlKokBfDgb+a2fa0rGjibXt4Ix
LW8VXpywW1Dtf6cKaIHzM9KJ7Uh3avkFhkb+Dsz7Evv6V2U9sNykS8imLU6yjojGADm2LuE/Heu4
wdBgHO+eukTXMvJZhAgPXZKrj0U7G6zd6AXzDVTolZHcdmX7Ik8/d2PauGDtwvgxUB7uBkwmKaL+
9gbUkjD6y6CrMr6GNHvIP3DHgQ7rhHDKDmIJ6S4lEIU/rBFD7KwdwHwRsadW8ZoRjQvuNDiGYoV1
YkhJp/igaxTje/S2P/UHIbQix8OmXrGrOfUnln4Qu87zMwRIKA1xvwtppjK4ukBLWvt2YMfIJVGF
EzpPxEM5jrrjZD4mXsyGFfOsOh4PDttk1WYsgNUwQIA/kfEy1SrnA7GFwW0I//Y1xKAs7gSOp3Bv
xEr2YQ++h7iOcF5xJcfZisTI/xHR0Spt+0WHWInZ0wl+AeJWg1MUyhBbst68oJm547cpuHO89SYM
ScDRg//uaeLfh42sWEEm0zICa7b0olUBcaGuEIY0TYuncRBXl4k/0R3TQ+Ob1sgpQ2NLWbqPzRx2
MvPnG8rlf6l5Iz3mvcZtSt6+iESwu1Dpmk++TTk8SQ+2Ic/u9aKCr8A7rhCZSt8on5s+vrsVsjnh
bfIb1I0Lr7tFgB9+zkXstUXBHoCpmw+cofN/9fYQL9Eqajp4nrvz6boeh1vX2sJRAu06zIQaWE7Z
BVAXMVnlJIfcwk0QrFc7JOTAbPX0u9kKLCXp+Anqw4IkyZj0eTmRQxzzvnEYUYXXSSIw+sp1uFb9
QEplsuurRwZ+qOdFE9SMLy2iTltE+5vXU16EG8y9n590VW0N8kxEXYM22cMagzEM6QHCyFqQUJiM
E+8ILrh6npPO/sXPhvW/ytB1tSpRDUVVQ1lvwsTNHouOI598IgyukR/W9lLQVLMMnVVSa5l5A1MN
DiXuKn5/EnXIE4f/T5v9+yJ2xtvoW+S0/rClJduFwHyvOQ3w9FrHfHChrqiLLEP/WLmbMpvjsyIF
73y1TknXEJm8ozg6ycaxGlCUokdnPMHf6XnTq2EKJo1vrxWMLGhIbdtLWj6sA2VhbA1l5LtvRVSN
GAN99w03ufOz+t10OVSieDzu6iF1Ale6rJqbI3Z7XSmcAf1cmSeHbMBX3OYqHXfuPpeKj/OH8+r3
HEr95icGJx7FeT4IhF9Ihd/6TQgoou6wA6IYDZ01NFkvijEXv5Im7MkRQsycYAcOXiN/54mQlEGQ
/wYijTospEyaqIqUS1mwYfth5n7iaWWR9IuqYjrt7rEcVNhnBs4OJahD0xoAGtL8BHwE24r92ydb
AVgBgUMFDJZQZIHpqYmkAOWu2fEZEKLtV+J37Hq9RArUITxP3CXjxKRr7VCHZKX23xbj0yI9kAx/
xf0PpMDbK7UQ2cC8PmXMimkGMsaluJOr86WGIohNkVzfVoEpXat5frENCTB0IDOFITGCd0R7I/K/
LLRWtm+9w9qQajgR/LCGmIspgZyVyckJcH7s8AUAUnUktfFdjB/CpZSKqfW15R7KYm+EI4kby2UL
VBhLGpiEpri+jk7qWz7rjAittGeBE8UJEx79V5xCLdhq816dsLm55MA+OLIQlLB6EhB0QcMN3uc/
SH9Glg36G1PRWc66AwVAfX6CaGarkRRvPJLlpzml60MKC1oP4mz1IIF00kGYnqj/nefXZ59IcfTE
h8Y79snuxtyf3MCn1Gm0w5Sve/2AtrvmlgGtLJn3u8u6QUW5xW4/FrtKDTMu9b2o/cf9d7yV2BVT
itSLPoveB20aQevxq8vZ1DOTLwoM+FmYwe8fcRcQT5sFpY6y3fEpZ0ZrHc6ty1t3zDjhSjzjD35s
rT2Zip2vPFQ9qsUbr7fzwvXt5Jnm+HWF7q2YJGvg2LP7qYhQpe/mEGPXJWJiB3VKkjAnuU615dSy
KDTfjSWgA9ElYKPfHCpaKyy42+tWyI48sJK/wR/BeUGuPr9+qmgTO46bFPZqVCZN1G6YwZBOVI7S
QWioR5IvyDHEfg0kazjZln9AK9aPT/GEvxXEBIVmzI679gDUQ4ZvPGmfypxtsoJufTsTsZZfMSQh
ZNZB7FTItMdtESeZ6vWE/VFPPgMwNZxxca/JRmJamHyYHITu+qu7V2zHyTnbW4u6u1O2t/cqyIrj
p/EYDyR6lWt5Dmlww1mN852ndnd5uluF9Cd0WNssFD9HHIq4yHWK4CuG+bexODzPBmY431vShJNg
586VXzADymVbxawDyL93OrKbd7VXKclZekKyTX5pyJFQtKnSBpKD0BCg7m8te1lyWZYqcmye6o+B
MVEcptvKjlxJ073t3CGN7QT9RSIKxqS5LHHIZ6DUJ7O9WgjbBNH6K7cqOPT6i3P/Qb0iEl4zWcx7
fvsM3EgAZuhESiYco5TM61ppeXG+oOKuVvdeYorzx1gTHDd4RxeFoHJmcqxTdYGVtO4fgksmrFB8
4HUjyYhK5WTYfcEvm6WPmJDM2UG3thIpzsTMHg6WkJb5ocmQVPvXmjWXHD95A7C0HTm99rXxH6Lz
ande2IMgP3XiVduR/FCUlV5pR/mGu5p6Y517w9QSMrb0Jlpoz43c1UHUUiJnLiRYAfn6HqmNGW5O
LFf/eqXh7QzK27ipD4wCu6m2wg3aVGJtKl2DmIOG+2vKKgM0GjMGSSz59mK26Z+si78aug25ITRy
9jzGHZAsNybhqqRvAI7lh1uI/tWb8bS6TOTTHUcaPaJzhLpG+Rt53en+k4fM1fgajLQuqxgdq2za
xrRTfYHEyaAkUQn3/vPVnRXq0mUMhbBljB4OUXTYkkF7fTsn+MPEUWeDDoXvr0sxVIGZbTiFgWoq
M2Mj03js5w8x3/Wr1/Od1bZby7gQCQhrMD0amoOf45eQfWCmXCWueX3giIqcxlSnqN5qwfu9DhVd
9Bhiv/fN0OMoBpUo9yyo8xPjUxvRz3eD7AQVclViAq4PXdkeC9w7+Y4znkqJgInBfW4NyO/RyaBL
3Os70oaxq0DA7lwaz0FK3sRERakUNIWCBwq5leBt0Doooj2LFa9xQbcDK932zZxwdGROOMy2yG3G
KNinoUI3V1h/0zcAThkdPrLug5H0/tPK7DahTfmYfsYtpugB2I6TO9PyOV7AdxTys5flO0zxELwZ
/6sz7Y75jX+Tv2Vv8xbLzKGNNR+WDCs9X7DJXk4fYwZyzHNE+2KXQkpok87IutbTWqXXm4oyVFxy
Lh1A32GCrfUIIMj5NnTG9u08cQHWt7Y8BUEw4qf2tueObefLG+AKMSISKH/pcqYNfHcwwmRJBPFw
tZpZDQ+LcubplXitTkrl1GfdFdoXcelhRtFbuv46coR3f2IZNkLf9saW31c+0LtyBnq+qg5G3t7K
1tM1R2X3nQ6WXk4yiDah/Z07Sw7DhjaDshIq/+TCcIaJ0mBcD0HFBTenp5Ay5TZeH2S1EqXZVSES
uIY3X+xKKCTsYv3EZcSyh3nfjGA47VcUqprkmu14PDXCWVJ54urUt2y2+CnzAdsmdiM1pa53mkpw
cpqJ5DAssd2haZBFI6e7kgecjNOMdAo3zRlxyFjekcoDtr6wphhfwVXL0jEl50ae4abR9Azdux+I
ipSrMhVDonXg3/C6qBG4/u+Plfa3Bl4r1dy7n3vyvX4JrQvpGOWJSgZcnQ+czaBL1zgOpZwMXRBV
7m2SydLnse1i7EasmqWhzo8nym/glbS/fG5sRD9auUMgYrLBZEyoxgzY9eLoR1f8RertEQ+0CEky
4PxpT9j3XIsvPu5NjySBGGUPe3ykNu7f2xTuEkR7ZsR0MthZ2QjyDf6acXncm8cdQcUFodzL1qFS
L7QGbzHIU0ac8AfYK598TNsxcSv9dibB9hRRvrHJaliXiF5ps9GtO3tBHRT+xlvGBa09wFilsijC
uCpVf2f74bp3aWlLnEcPaMFMTXxBshH9VDdqpurgmfW1ObIHSVDrPJbiuCJP64E7RWYvAUxKi6o4
4RurGp6T9gBaD95vlrx41JQuKWCgb5KkwcMyV7Uy0YClMDzkhO1lAKg8r9B+xb+21XHarKUEopja
oCTSjNKG6qv+UOqwlgLmH4zi6BmWbEgN7tCRsy67zwYUKPa/IY5QbBb2z3ppPEmPiJwzY9jeS23a
DcMsot5BgyxPZhXrATHHN5pNRPvvwAvF+OqgarxbFrdXwlZuCXIAGIGFsyu3SCtTrdXz70NsTqSv
kS0Hy1VL1nKcHWn2sh0iKzFLzt5zxcCqlrosOyLEIbSmhRRAPEDLIsEiUNHybDRqKxody3AKGmi4
3gcqvP15KsEVVPz0cO1WqUs//JJDRNJavSvyVRvnsZRNi8IB1KGDyCSO9V7SnekBuAwzYCEpfxCt
ecVe30ppjAmkp/YoblVDc0WK6zLFeu7IRdOmQq27N0uFIRTxoXOxX/FisbHYlDnG32JiExaMgrL7
Agaij3KT3kHIzwE5LUBfhfxEvBcLDqoiabu/qf1wAVyYlCYN2uiEthDVVQxkDNMrJj1b0xlSSqAW
zZkM/caSUtRykMVMfdoI4ehz54jzROZuFBWgHQkousdJMGJm7oq45FjRHivnaYhjDju0tWi5i7Pj
Ra6vIaud/7wd6FxwYUc3cd6qqvGafvET85mOAnmqu3QnUxXPPhqdVaHWTO/yx649aA40ZGj4rojL
eMiOmVi/NSXHqCeKmXqOmSnSzkAdcwfaiATff67HQxAs0VMGTYfEqKbwOr0EV8Kd7wrxZ4BURJUu
G6wikOanoGHYi+ZcY+jd8FmQ1ClSQcH55xC706kXilbmLEO6TpsnZfqfkRPcVNIRPXkMYCetA+UH
Etqz9TdORQNLdBRbGVK+IZDZriCs61ScE4aRW7fE6DfwFvEvs035yHdIbXyB2VZuipqtt6YZ/WGP
j7oiaB6ap8E5EOOg8wkb9WzlDDhK1c02BysBwQGRpM4nm4f7qGTexUxKaY6hbxzEnpJgTyqAx4R7
UEU5SaLKWx5S30CvyZAfqCU64F7tvTiq8rJcKqReWlFOmzq4Tu5/VvCXbtSojCPepJmzC6utiqHs
YKS0ZAD0jx7XVuqakrSVjAAvXU+rNG46lWgwTAfaIqEmopxdSmxJtdRb8SW4afNeVfneB/LqZKhu
wfiKwaMY/TAETcvdicEL7C9+a03+ldByDjh2HRt+eH3dCJGHjPgOz2GoTwGGbnW1F6uSh1agzoFY
ygkOrXHFIW47bcR7PUZzZ/2ZztqSfBnGfS9+sI57+rnmd+JXiH5ATS9hq+7rLH8gMW20HtVM1XUu
c6fWbVc7OjYOVz6JlNjaFwdrU7Pn5vwv9xt4qJ4EZyw24/kTLWukxanvxsZXJOIPSJEtWlMb4AmD
1swDh9VgDKvEgJIDoWNDFI5JQ35vEJPz6B9irtNhZVPxOIKzDxSNn649nppjpTKnmyR9MM4fUlY+
63u0my4gIQ5A7GcB3NzJchZmN6QOJlu5at++wFafOhOxtezjIfLlIfQrbDuxyyf3WehGkpJO3xWw
RywPIC5Ce3wVjOKSNywxYxvCEbDwYjginS70qxJ2bt4VcqR4Vl5aviyfPGVeZDUVOlXh+e8qVhJa
VjbWBjgAsPRM8atssma1etNffoFNacmNqpQL9AyftkzUEhUIBXTQEPoZGV2xnTeQ8MKoo7gmUMBA
+HTE2I/nlLoE4uibVWJLYZ5EXTQ6MByn+ryAMhScRzx9Yx7wMfz8RlMvmyE9HF4mi5rnpUgUY4JP
03Lwb4HuWddMI3cBRToVOWOVIIuFwsEbGkyS3HlAYlh/AOLLrBdhBKudsNtNk+cEcMKfUn8PmmJD
qfAIHcLDoDffG3th01nW2hUFu2CBEdrza+Slv6c6Wu5+kCwu/ZL26RrRszIq7avH7nzil0DqwoRi
xI06FLPxAQC9HJWaimeMyPRhYTO5Hex/XdVUd68oA6T6LX9R5L2yY+qePf0WhKq1F72T4NS6h5Zo
DuLTplYUvluA5xPmnFApDFHBKKFMgwMZ6uCtzo6jcDX01W+2n0f0qIJ8F33pGuI+sph3TqTanyI5
h3kDlg/mhrDxWM+l6+IFnwADUQl2xKxGayaWQhtCfg0BzC80Ro/sgwOooli3rlz5Zi62DAuWiHI1
i+Sa97cPNfEM2yJ8OEtLWnAcTYrwmM7UjeXqHyeHQiVsdHtF9Vrh+KmAZGPOCYRpTXd1YNSNZpEx
vlgcxdtJzfPrGukekUibgrVoio5SLJJsuj8e/VqRG/2WaER3tH4xsmQyf4mkr52O6IiYGex6RnfY
HfinYTqjg0Ar1LtfA6KhMwEGJR2s9JoIhMF4gLPHGxSdcnRBhvQf7lPycVIbscGYex0zd0i8OCQn
wcJ2V1zHNTwCe2fGuimHLaegfdw2tBzEIJgI2yEFRqTCebWkR6vVwdRu7SLWlStHiU7qPnFk6uH9
ykHzUoPRsLDZk74JQx4x+e/an5eoj/ba165/d4NUHpzli1i+nZBFts0JR0jq2xZhJCluRXvVUpW2
48krRXEQ+PjwOW2ZdAjBbMAqELgap9KfQkhXaSzk9DyHZQ/ZXYpfPE73wz/tz6f5Bkw/Q5YS7DNH
pdh+Q4W1B/Nc2BtuvMgThsHzStmM9C8UQjm8gf/+hxN2hS/dyWe5eo0wTOJiYAap6zxF4P0eeyDK
vHE7laU94dvif3Q+PkI3yeiIaPIRDgvrlgp8ggaDCokoyOcUl95bh33CyI9qpGjryo2TOKPLBExZ
+g25U+Nztv6bdgWexQhjT+nOOTA7y1kIDGYK1A8R8ryGOLmavdGbumMJFNOQos6rg+eR1wIZEPj4
tRaO+vZMC0V1lNnkP1ujuD4i1BooDIeOjhF4KVBmxsmCJYeeVMr+y5K41Lw+3v4LbWuxPawP/CXc
LJdoV4S5AueNgmxGAQRSdkJqozs9SiJp9D+dh5Gzsr9UI4fRgMIz8GMqVtZx0SPZSCTK55MKQmUz
hOag3+dR/P6HjNo1sQW24W6Ysrz+bkCBzD7FN3o1vjAmHLrmaqlrI3FO/IrlNl1CGBuJ/FRaaUAU
XS1IKzen4IA5b18JWBJFbsIEgFq9ppobPH9C3EARuQcJKxHtwqZiMMUVJvZr/20Sq+fubZQSNJ1v
ZFLNAN7fXXIZCSnXIaFhmjTqo0qRUDHKeBqL6lnWIIi7AQse1eFvQLpEAmAiMtPRNqee56vQRvD1
eNWQJOlPSFq22itQQETeXxJCC3y6nc7hB/+W2V7lOgsUaxh7swdSTu0fLp2NOeH3SlGRreVlqDkm
1CJO3cfd6bWbnhpBJzvAmeTUpKqKMM9cUHTTXjFTdA+kPcB4gt47rtjjDsL/IAsMl0eyvJepvvw3
oDepzLnTcHlUXLFp57Na/Wd7/WzN2uRa/hYT1Sc6txU2FgyDWM6SzWxczjCEYY/IylIQ/H567d9R
tmB7oMzGzOlEUfz15xMSI5gsnP46X9YEEKSjzo80VwGpXNNTyGbnILmmthtHePPVpE7P8sF91E28
6NfGB8DOy6nFEYQG4xpaUtPYgZDuZNCcNR11CQZvlTGwrTwyVDl1iEZPuUXW1JreTaItO3pECbDQ
DiY4oK9GxhsvJTm5EsVadKGrFUZwUvuHxCMJTjBVYCRRKk5mt1kP4Nnko5NFaPB7d7V6QgT4ktQz
kd2JducJn5yrOgOUFeEj18ZIMRh+e7UnqddL1OcILC/xYGCXsqZubD9UbMnYx83Kzgtw/SEmfSdv
faGsdwtgef80UeNX8VCJYgdla0gKTMJCjDLWpD3e90bT9LhS7OdhCm57WsliUDoY01YPQYQsKIHD
tgmXhb8j6Kks1D3AaHElzIJGNlY+IYERUMlqWAxmiDI3ob7Fon/h/6INdtMSW0ZOKL8gB+3xuUWp
42D0hVSwELnrQPHAsW/ZvT2zWgrwCNvpqifESmHatoyOn/gh703qvYtYrQLD1SnoEdBKc5HhmJh0
JrYQHBhuoOwqeqMY/v/hwnq+bxNUtCx5ZatZlJFPP9JguGZpEsVEb04f/hT1TgFggKjcfDogmf/M
ds5//0OV1ZzsIdNHMmUSskigQIXiYVmtZI2jFSXPNRcd9lfxm06grO+M4X5Y1QHgms9WYei/yh2t
sdl2XaW22niQP6f31KcY2PYE40/O3bNeGYAapswCYLGuwR1K2K27C7FG3X4M5kaNzgGrBUaq1DvQ
uR8MCDlbMKdCQUaM952IFg5kfG50tZK6zT7j0tx6NrF0OTkHZoW34edTQNhCGRE2ykVmJWnBD2FL
RRfdVuYCsxOd3YhkP2cHXgloO1Qupo+A7U7+uqjjjSsqfh2xDcJC5MeJiBDG6WGeBtFNXQ+fiFyq
uM/f3JO1PS0/Zn4ucgvNsfQfnBKcK2ytZ194gTxeMyfECZetClIdHqWWGKf1ltNiSQR7NNl1ydch
WrvwtEAekzg1OrP0qM3OWlwkvmdMxZJl81r49ayYzp1tz2aH/TI2kc9xPWHbztHfnXhDNZ0U11Tn
UsXyzj6+LzbYZQ0yfY9PLiGJXpbJUESqvwlK5CmclQP3J2eT5O49Ya38GcIWyqm17y30ZQ/QElo5
Lfhac9s7lB0rSrOTZbcSs6pTGr17KiQPza72gMClwt2M10f6QXGqHL/joHuVaBKC9+hpNwr/Ib7I
BndiPenWos5FVmo4d4Gf7XNEtT2NlHSSPrpKr3iAl/v/utJIl5nqFls2a7KXXOyH9EQMAQzzDt77
zNTAuRfminLwTwuVi+Jqh0nwAcGpWctzdUlHFxTzk/qS8DR/PiowehzChkoRIeex199HDRowExKa
vkKd5/ag/13wDzbElFmg4QqTSkl5wdpyTBK+Q9AYrZNrIs1HAzcE+gpGkpA+o4HdylNBZncBNDL1
qm0t8GtYbKhlXAsO0xl2iH0XpS6wXeoFKQiS7k93S8KYpJUd9f1+HTD9yUIbgMAl96citpeLA0ev
ezTw1w09TgU62IoGZzfMvEAQNutj448pQ/YIaRrOiP/rukPxbaFYwLAJ06hsrdSk7XYVhJB1vERD
wUb3SQSbt3+3TFkvXT2xNOrONGcVAJPowEb4Dd+oveoWEg8Jk+lq3/3tSxr4OnobR8sBAgZJq5EP
2BD8MB8Rf16YVoxPjZpLsYdMt3sufvRxEXiv+swHeTFtaxjz4jbO6CcJEYpcCEvPxh3/WIfA6U0X
79QkPBpzctBpS5nzLOqSQpyIgimZHTrSpir40Ta9HWzX9b4SFHCaoL4C+VMvkO+BKvntJLH3Wjdm
/HPCUWe1VIA1EeCOkXqueeTby6SvRsNHhXWlZk0WPjENKMwpFWbiAXDWvAzRwq8R3KCpngkwBmC0
D6iclyB8L4ZmzCQFnNZowOODcO8ySVF/aF1qT4ejrS/yXOR3gV92SHOm5J+VSDEgaiAAk+mK9F1i
xvRzTeVbXdl9HFIxT+Lf9NZJi8ktU64Gj14xy9iUEekK6R76d/gGRIzUrjJGStjQ8EyCoyANkfq3
gmHoeU2byQI4W/K8yFdbdGvMdCuczM3lGmmGkLEliSyEOkjpD6Tfah2zf8FSBqbcSuDYYCJR8rH9
ppNC6zmuvIIfP3p4CZ/napHF/z721DxYgafmEJFRT+dvNh7uq7TOXWHTf2ogdXu1E/E25udmFUPB
C7BuSoG7Rv1MlFMOhB6SWaby1cS/eURUfaA9jtcd1jaC80eqjSELe4JOz92azOvSIFH08aOjwaXN
We3y9/HOlFs9j0++IqOs19JJXls3hPl3IpPKHOeH3d+tm3sxqJnrfHGXDAjQmi7Ne8fxkxEX2Ehq
L4bSYU8E7+QgxVYgVxbU+mIdwUgjnuN9rySFYrv+aaSFLcCqqeWIlQHz7GuS5FgcWjD/kJc8F6mK
sg3tvZNxdOTjW7dMfYjPoYaT+rvHkD0BkjHeOeIx1RkeMRPOK/btMd/0QITWFSdcxJDbp+dRaoOq
U5H1+k9Of0dD5wxuVsXzYfZvcFGTGe/cPRdmMGh0JiyMVMo/vbIl64mZdEn++QR57kI6Zq1vlryB
nRwr1L4QvJBxGPiGsTMXTukuny0+VxgxfKLMx/WJBlsiTxH6BphrG351IXjN5QPStt0Paz19vPK8
0lWzQK5iwLsl4mbt1Iv4U37u9zPquJoog964h49OxY6U4SbGeMx5avbfK0ryYhEmS+2gv4bilvwJ
yNVpHIxE9vIdkk0FmQk3XRUMAE10GDr7QieZqRNE8SFBL/vxYazdMh7l7MAbV0Bs9D8xOu2rNKzy
tPrH3GycazGR8vem+CziZrQTtivEHUd4WrOUgaXPb3lKTnLlrE4XEoiyGGAyvpv99TvojxnoHovL
f+VjpK76eIJ1xt8WC/rH1tR9lLZsKrUIBmcVKXXcSyCippxY3OnNRnalOu7FAmIDrjncluhuuUkM
AgYLNAqto1803t9m6hkhQdwJeQW/k7PQldzbc2ZHObvgzCtmZyXY1JakoyKjiSCCsj1+bZywXKiD
LInDQIB8koRBisIg/2JRRCNtR9TxG0Xv4cqgA+Dh4VMx8f3IsPtcZ3aGpurlnAVOm6gSiqbwpSM+
hPyA+CF/rLjjUhPK31nmkN8mMTp056sdlvaQFyFRAosc3TzLyG2Ijha5jX1lTNcv9otjOHUpI81N
ciw+nd5doL6Z9i/rUyGLpDpddRblrPiQJi6NaMYoNhC8Q5nfi+e48lByDn7oqx1FNIjleBuiz6JD
nA5cN/GirZNTr3gasGOgYtXKXF5g2laT5WmVZ8m9D75o2V0GaT3iHKXJK/pX3+ov3pDaAaxURiBs
/GPJwHgzQNOrcXgnfDqbkRPN8PVJhJienWGRBJTwwGtBTFrnkxJLGvRdxuo6xS1gRjhPba1urP8W
+Niu9GZZU4to2I0GzJVRZrqk3UiPzzmy5yu4182+Gk1pA+5kT7MjBIj0SytaRdB0FzHDttb/AXGw
q7ul+QFGPvMnyWhoItaW0dNr5gsSpGESBsMLwtqb796swlnGVFrhcRfWW1EWfr/ziM9qqb8Ehzia
niTTFv0dOvPr55vWpeCpWA3dRVSyYJePzST2U3ysOMsOy8oh+OU4Ei3ZMe2CXeUMu6I00FdPhrC4
csPy3ctQ3wGnydx5OvrhkQoj719m8ZALIaGZVsCVv/118Z0rD+N6pH9FOfRqWAC5xxXsgIFU+qlZ
MNpe3OUc06ksGVt1RDYGzhvDMX//ZQ72UXex6tGj59wZq6UA3Z48gW8ZdDxzuKSGdAtjxcmLgRtv
PoXhIyEAAMebWMlNhy2kIagjgVNjChUOTeZsbVw7adKI77E+6O+1RBpCcLsnSJDvZYFzuVnqnBTM
uybGBZFSVJg31og11hey+S2qC/eEChaqHD/8dlCMlPE5WZneKY/ZHifcuXCfpBgllf+ozQcjcRj2
z+/lozAznSZLmRcCKM3/cPrYrvX/vRLHK2/o9NdZ5FZIUTObZFl04qngNC1zOqaezySxBDZCWe8/
3H0znSXwXeMlTPDYdUTaPL/OvdWi+WqQxlykoasHBFG2dj7KFTa9QlPOnW6D/B/FV+tZky3bqjsT
nLi9SqTOTfMQTCyv6OGBKQPnsjWER/hgU/BRv9z9IIj0UkDs08Hje9A3IXBi4XUG9GU5alU3BHdv
MEbhnxpvyAw2rypWGHk0QTThYL3uHvcu8XZ9SQTvabuTuIrYdPeCl1QOyGA3i3rbq0I24OBeVK8G
vQ8ur8c5pyJDoSUBfd4O5J2klc5jX/0xUwzjmbKAFCjhXH3Qi7kqwduexFJcWutgIX0XYAjjTlqS
rQBshqPve20HtDGgzyYBc6hkdwTIDHl1eXNeYBU0EKCFn/Lskks/1WiiEH5hoGY/0IZGshZLxhne
h2nLXTppzvTvJmY18Gsb9LDuZbduYyx0F5i8l63Y7q0yBMUHde7hyC1oUF45GS5Ffx9FvSfkNOaf
cz363vl1RHwjtfSLIPyAYpGI2XPcfnar2Xpnu6k/5YT+TjknUuVeKHmmeHxHZWtymD+jju52neyD
4eoxByAbGRVrVMl+GOorHnSgBOm34uOnXieh9bzKNtnGtOw5VRNz27nJf//SM/UE0EQItiIuLGZs
2I5sPVYFaXgvrwMI289wmY72THisQQzaAl/y6T55a9dDkn+QUYsdUIr0lc4+DAlnMRgEiBmBcf+0
AqQ4G5TN5IyzhJpJ5j+XM/4s5kgHdBfdoyq1yYu+qItWwl3j4zTrnP9+yybT7Shefp5WGVmRLOGu
xocManbvhjnzqkmfRUpQp2wKPYuCDn+6Nns8Qk2IsOW1L1vGJMlsnjkziL9/wAIdh6ccq3UotLMp
0Ic8Se2TCaw2qZvxl2vUUWvlHmz22fhL0/b0E7ryUeFm6OOLVInFsA6PwzJ7LkrGwPpaJaqGIaZ0
yMir1thltjTgPH6u9LrI2TOeo8r9SdQzZ1V44Ls+sup5KIfKVHqujC5+NjtBENFQsgrz/m0SiYoc
2Z6XIReaOwelLOd+hsWxFKQxUtfRc/PA2/zNpNPLO3dRpHcp8qrR2QjesJKsPg5OES7YhyPwGwOp
GFNCcLt7wwuBJvpy1YDi2RRkgwZwQmClCY9QgsjduPKaby5/KfQVE3l50wnD6sbH2+U902cn/t0c
mx2vzTuRN/ggCyTb+p/ypmuOMD26gR44Sj82/RQDhANXJWVE+WWQ7vHUSGUqxynTlaQKoc1v4mZN
T0JSiI3Qe7WQs/s8XgaVAanZoEjVqOtfRyUfV7n3weD7D0AFju12ZpwcTmZCg2+ymGXecDlPUuHM
1luaewd9p0+5vXaoOctVbnN9xtlJ+0NfcelWugUQeqgTyxgoUBa/dg8PbM9IcS0T6uBixmTRf1M8
YGsXThfiV20sBAV881HQZU6mHlMuQuOY6Kti6bcW1CrR5t2yz9Q7AymlA6WWrLyD295H6QUeJftS
qoec/SVmz0zL3yy9z704k3b2JbfAQg+VQz6nwZi211rgT03W4mU3c9q1Tw76JTsegROCBlMBcU0E
QUp/9wWqiX2dIAxykhuRWOfLqx5ft8qwltLAVJPPLS9NTfgCD4FwBK8lpcm2mz92Ysrb9dMgrqmP
MvC/weMwIKR7/6axuKhp1F7NZi1NsOjNqNedylHeJ+49ilCEcdMrUyggRxexBTeq1VpC0KMGL6ac
oAhi4Y7s8UI6JJOZ6niiosvE0usheC1u5AQHE8XojBHpduUCDlEFxcKF6IhKU2ZyBqhVxzhQItCV
1jbF+ck2cz+pktzEP6QNpXkzEGfkFVLxI1AEr+mRbwIoCMQxVaF9WRCiA39iYPFN+Qd3DllWUsgU
XIpfgrPHdlvjziYqDSv8i79PfiwxrD5EexqUAUXnMsdlKC5iK3fatiSgVOzgJR8YvZ5lWbK0Adoo
iVy7G5JtkRxBsGjPIBGMbAwYZkSpbTUTqcnJd8W+p15qSVMcAMn6kqWCAKX2J4KnjETsYukPCppg
+uKo/BMJJj7Z7UGm0nqe30QIHIQJiO+8HfUOp6/2cPJ6/tDAHeYWhus4u1vMViVQugcF88wxktcX
6OSHAPRPd27co0oUdpIuIewYsu56v4f+0y/g/V5TpLie7kXPu4jJsyyVwuSn8IzuZa9hozHT1ptR
7RSGs6queA1HSgmX6WTaSeJpoeCfzLLUZP5/6nXvCs159bBr4lync34K/q5+qU/nkWY62bNk+R74
tBsdb2NknmzXLhbCq0Q1JREd8YFg73tP6WGPe4HAgC9wttTcnOJrUI0tdKHk6Ts2gxWKYov+Olof
nt6sXsCfhe3w8HpuNOniCSfmZ/bIvTGclz8OBNuvXR8iwI4d+ORip+M4e9QhcqBwNwXkRUYGGUPA
aAPiYofiTVkp9VRbwjcpwtSHua5ZQ72CoJS8SRe97fp7ceQrVvQtJwb5h7n0mLfzqWNbmHQyvznY
Ix0Q6yZD4CYspAbHJ0urPSWybL3KdU/VHhQX/BB6CVezIs2DNHNpcDrkzCqD13U8biEtxbL1+gvQ
1w7fA1BbJKWILRYXNOipFULAOGTFly+0FgFb5Fts6cwq/4Iw+nJchjDRner5MDu+QZUQ9saqHn2n
cJIuNH4ufLoVN/PTcrdoiRJHPAGYBJ16ZMSwVF0R2vbzKoLMRMHrMJGMzAa4+ONEZmDMn6jxQZ3c
pGYb/RqmbaVcoALOJ8Y+vTC11krTYCDdSykcaLX9aHmw4aYEaAfcgTwtXDgGpVj+rnLHBiZVv4E8
M/UvthWWWnVYlMxeZJ8iqhQcyo+nfCAWyafxObuaZf7UKG+Ndq6JZ1PeTxOKOL8MW/u88jMFqrD2
2XaKdv2Ea/QswuCTW0d7tTMdZY2oXkp+KOV2HKPEyZWHlFtfl+acvyplYXhmYLScSD/hb4pGbkn3
3Vm5SI2wlOgR7GZ0+3FhiqiEk82XsaVqLnwaDUYk/fKbTFYT7o9LCdEfQgFlX7hPQn7L7QuNKZB/
3hTymZ4F6wkBO0/9XruDO4Q3Er0pIPn6opkHbNy4CleC1wjKOdVs3qGl4uIjVyJWXLGlTySblUTq
NPI1TeOx0eRSE+MwtYqWiVd8C+vWjkvD1EJTcjF9Frg10hFJcs/Tp/kVloqOP51RcblRbP2jfxS+
9zKp68Kj3NSP+nUvgvj5fRiIl93ar8nlKIf5RmNLP8UvIR3Knod4R0XexK+W0uRDbl3C6c2ifFkF
obYEu8tFi0bTVtZw9+F9MkXXlGw5Qe5SpHsl2fi79K5OWgF5TrofiVO/a0IzrLA6kiFvZajnj85J
kcSQrpWELt8advVmnBHLGlotDfnJ20gZU3FGS5+d30GetRahXq0bH0q0W/Gu4CsqR9Q6U0zbMV75
C71CzhHZ6sCEXA72RvrAIU7Swuz4jBKUGXXfUIm/bLoynI2OyZUGEWiMY9+7jYQH9Ha9VL4LZGER
/zHgR1NIBJLWAtSecVPEZiCjfoA0s8rHBwxZit3aLpjnebEzsqlBcUd2rqh37xbg6VRznq7ppbEj
8pG1tBAkGs3GfrX5tKWw27TFtcuO83JIZStJUA0pJ6Sq4qubIs8FWJPqy8mISpSMSdVPqsFvGEx+
Vrp1Vxgl2vWcr5/VKK3jswEzP7LSQua2vYEQ7do0CwxiXVlXMCsUl8gbC57e5xvtOELpNryT+bti
7tyuCRELcoQFgI0bqv8OLkRzQqbqsTjFWMB/1kZBv+rJKcDJLCwTdZiNo22aGAWg4ZW29up4CT8O
rXUBBOvLRFTNu9w8eLDV0kVuVEI+eu3JmUgXFY0AONA6h0FMPKmHiY/nhz++eM84Q8gWOfQYWAMW
QQBpPQhyfpmN0c8MsWXkaKOp9QwYL1Hf5q0b7p8z7MFVCmS/E4WS4hEsWCQmlDIdp+98cjlVCCXr
sDIrB7tzwUPYa0GHi3vawljQXFBdxhuQlx+UZ2NZgDkW8fqdCplP0gxDfp9hykN0Cw812tX3aQ2i
UBe0ERh+xH+zfYNUjCl/0EGR8bgf/9blMffHHQOJ6X4prYDbGGXT4XMVImznH+i5MsEwctXKJiYC
6Q0uvK/BDxEXXoRCyEeO1Syl1guqdWfdzmkGRVRMc32aRav5in7qk0R9E2JuyrvvbYv9eBFZVgx+
5peJQbj816Oq8d1fo/rW8pFYt6zhC0wDy9h2C6XhQ/CqxQY2CXsc25QM8z84QwTbRq3lSinsRCG0
0DkA7LpNvF6NQvHPt9tUyhj1oNdVh20CkFft9ILSkAtpBZIEc1sIj8e81+8+cXGukuSpmV0lTYlx
4TIvh8/+SHbIZa6LegAUVoCxEYdAVRW97WTARbt7IkZgk4C4P/sbuzrnxbcXl9pZt+kxV3IGexTj
ths+3+JGOTRsNTE+Lzoq1A2VVquXHqL28gHIYOJzZsInBr+D1UXUoJ3jUgODRkKVFfKgk/B60xf5
di4IuSeWVhDXa0bHIYL8hFMem0Icd4efVbdL0+TCGxqsbUc6/8ZLOjHKPQF67cGKAWRH3FL7deGl
yoXZfSPpZnBaC+Vhsi9mK9n+bjqs6bXJ32NmutsFFTOC/PWYJscYP9V8kEnA8v9FNd3NrKeO0mMp
3uJIJvigUO+e1GbJDbSezRif4CQFvMhiDHnTE1Ec8KIKl5o0OcBywcHepvLoLbvk4IzpvZ/kcsA1
ff/OXE+iKwfDhNieiML5M4J05kS/7FFZRFPYLNXvnYMmwQaQd+SoHCjftOYdG4KnhcIk/UrMURCW
kzEFaxY1iij4swc4YFM+88Gq2nrSGeme+gXSHZw+xnPRTLztxxP9u15OiQprPoDXrL+3vpu3Nqcx
KWKGnJbwZxSx7GMpEFOYOuAXrDlSheiZyymlICb7pSwaRgos6e0IFXg3kCaEi2WdXW8D9jhnhziO
/bKi855m1OxAbJ4JG96I673r9UDGJ1FIu3QWrKBDU82QQXnjWgr+A9dWUU75no817XuFaX3oe0jp
TizJ0YLlGwKl8EuU+mL8VCI6v/BfkThJ9brPApdTpJZQW5Fli1Z9l2Nc4wJr1pavBTCg0+ufcNJp
lUBkVR5Q+u38EubQJvRqWd1dnGL/OX/lWwLvjW5qnblo7CHskTwuTJ1AmwDfhLLbe66vsvVbLe+j
xPxLwWfQWtdTsjZFTKKRJR2RUdOLXziCx0oKIP6rB27vx6KD46YBliWjAPvJX96jSncFa5mteTaN
VzcZLNr10aGyi9FO1hjXye+3nz9zb3APXxuzhP/c7MHJfnC3QDjoiW7dpzXlJ+8Wl3tv5qy7hC69
Zoc2xgmh1yCvZ+E8sAedD2kfC/FcowpMSQsDTVXypfRz9oQ7c5PQY9wrR+F4yQ1CI+qz43QN64J7
ApapX1cGDXXRvUGeSKnprwftXKk6hijtOvC040jXDULFKyO/5usaO1YYdSB/qcIpx/OM0EGnTCeg
/hqHXH5OQ31DPj1967GHwAHEjCvXOByHG1KbkiVDOjc3Dh4MVf5XvCODs4CoDYAur63PJw8KDTkq
IAHuplv1b2XSC8QgwNMfWCnpH5G+E7NYmkIHx7Vy6uMIK4CMasVMPtFLPgtlE3PMBOb5BuOSEbyG
xemuVcBMHwt0YMAkVZiBjMZ/aEL0vlboHYlxtfTj7PnwY/el8InHAtbWFUVWnCfJ8dn4aUwWDIB7
7zT5L/7m1WHFZN4CBfI09XM3UaYD2moW/yqx/D/0ZEf16tbOX9qsjbkzPMV/0jGN68xLndwE9DhT
CtMP/TyFkVIlB3aDMXUT8nsStw5fOSfF00dr69FJ5jrXvx2VZRKUx0Gzu5dkcYOl2VLX0c5GueiO
0lk/5GENyeuOUqArnq/ApIOARQPtApt9Ki33RkYFxakwiUL+ymsGSeNTK5/ZOAkY+fqYBYwgoREg
8fWmunaeYk4e4VxjOWa4+WXtCtJtKV6hj9UDuJr3Y3uFTFGtvblrdz+7e7a33EZJCxQiwY/eHLLV
ZNq9C0l/5YDhGY13OWUX39Wu1whFG/rfIeUVM/BCwEoddTnHr6CfYgbw61JDLEus4carr32GxYJp
l9QL5CUH6QZrTf0e4gLm/NKlN2FlV2ZPGeyeCDr8vzL/ZPGTSupJdnwtGsvvDATs+sOKvomRaqIA
1r9tJVMEbAAp413sM2ObtTOp0fr5NgLMD83/iY8D21KqiYELtQGCMRyqGPKwLRprIlT+NEIz5wrZ
SudDixKxKduWHeQQxQUh4ZNlrYznt6a+FBC8fgJi3fS2xs6jrMtZ92ahcz5nhV7J0Xe0GTvPWSJ3
JbDTT/Q7j0bGcLLFqOFl4ANfyX9ljdZ8/snqZ2RF2XytSfWF5aBx9FXWUUG6k/ZE/wVDKdlj7wMR
Rd+e0TAWZYxJgmAzlWHc2lWkhh8KEeuwKLLETkZqhnF0r87i8rdkKfG01DV28IB9tjel05AXViwT
cU5EVAn2we/JV46ux4YAvbEtZ1s3GdDFXAxs5eLjWMVtOxGY9+oO425DVAw8yaOP7NyOnICwCdRL
EOMzbXr0KEu14BbwctrnvvmgF3FVTf4PYJjJq34rJYIjpP1tvlE97l2cRQsCoy+ZrBy31LpQg4Cp
eUaU8vVISC5PMhwdfahCV7W1ikHmUR+i1GtulqRVqNZ4HDtS0t7lrSsdrhOF6SzHWHlNXDRg5B9i
IyYT+F7eOVB21N9tXAUoP4ArsRvtZfh1ACrulggYZ5VHrvHzidVYStOlHigI3Z3ylaNUonN4veha
XZslzD6jlTL11yoiU3lr9Ve/rupTV2FW9gLYH25hEXYhmqyUZcWXw5xcfc2cBPaESjFjuIHC894o
yJH2ItEk7OGOA1y35n/HrfOJfhgQbnaXgfV/wD66A6Q4FSTsvgpU/qdLQXB/g2lc2KMs9DR+T0Kg
9k/CLsbDgWGkYU+6T5AlzGbjgwc3sAXrOWBSkuPzmsbKYqXkMAA5eyYz2ytQYxhwDEZq2DKGQVUz
qoB4lkaAw6dcPm32LsqsK89ivVB8kwp3sObFxnVYo7WRy44960eVuEF8FVwWccrPzO9xpjY/8RgV
xyA6cdAIKJ8BMkv7IZsDoXdML7w3VGHGoUnn1HDLhgRSaP0TONRwkjZEuFwgTQlM6ZVOctZemjCo
WxGXvCCyQEyMJxkc2KwH6WQex6uu5z3cuzcBt/t9orpf6G6gi/kzZFe2T1e78yYRwVhi0MhNhqkL
3WdtA9VnQYpizTxPspx6Un6RYeB9JRYPyDyq6lwmVJl35S9uaOAMUk2dk216UBljaOPt5eKfLvNk
fGQdZ9F7vlgZOVATg51bcW1vid1imF51Ad57zPR8Sz1WJwfcApXmTePahcHnDOCbcEWDtonoTs7H
gFWYR/yQZki8U6ibw19/Oq2VQxIQIE0EVLhb47guHQ5BNbnMpOJTOhx1t3ow2E6fGWkkiK7fiTbY
O+smGn/a5u1d3Lf7F1uj1csqV9MAV30f33KX7pOyG66rfPQ5rpPpdTwFSfyZhVy9tpBssz6JbOhJ
dLRBcYo8l05+0Ovyr34beYs+9Y9pSBScKb/DEpxaLVQ4QZs+EigGO93YQ6WsEB676jnoMLbkcyJC
t5efdo3gaRJNbaObIF992P5ExLnChK/sl3dR+RFWlaFsK8Nab9SctTLK+QM7KEJeSx37pKpmkp9/
i4fUuDglSxGmvX86PdvYP8QlGmyDzi+CSB0kWiYkLr9V5CoJrI45uHs9pyBQ4owdnmXfO1fuDiD6
dLyRTIE8hvrTzMX4AT6JkGHY7BLunxzB9HEmHaN3O0FO+wyC1IJ93XLT0LtihWfbDvN2tCs2TnMW
o9BgirPg0VnIB+HEH7H4fQxqTVnIPN35OcRIgNuYnqzMvOLCPm3N6mi3F/KDNKszM4O4fTeDxvkC
gmjdJDNP4ivDFjg/YQzWR/v38M6Y+2O05V902nri90fa+xRYfKtQOhbFiVE/Rjo7xeQU/0Pi1J5N
TaFWDDAIXa4nFK04vfIFaonwaQn5lUhsJChs9iTKnXCUmMAZYRJY3Eo17jkQLIzPepaX5cuEZyLf
2LVRI9daEzsWadwIbUXHaSZYbETgxlYx7iXQ+DUO/rC0VMCMfJ+KicIQYMGOF1igvzyDFCKPizOc
yx2LKw2a3vDsnIQx9tbSVoO++WGg+6OfKpSxjn/QFkOesHeEvQ3KMc+DjmRBd91z5XRrhICFhkjS
DSUYjtA434WNsvwtKHaRVnFEl5Sybf0W/n6BRLlXFWOGCk0cb8Ccymodl0417GoC9bg6mN1fgmeH
GRyoJYlxPUbQMeXWaX0SVn8SWjq5H7U92elmgCNptD10H2wkXSI4UBdsAV4ymbiaaApOWY7wpYkR
LEDNaFVeLrhbNWZ5sj6/DUX1TyOqInS+XbvCUzEyrRGJT+0kHgFCjRXpGjpvDC+tokgY1de13+xo
omyFGnhUGvGNLGepT6feb0SvfeRpvVYjbUcoAbbCrsOGFsBOffvKjTh+6fOp09qV/Ma9VmWSZOBH
CXiMu+xOFrSevus+e7LfO7IYjhiTQ6Wij5KpAkljpp8hnRKtGMLcSPZuM2LF7HDFkWG7D70Hjscy
JSrqJu7Xf/ZvNnC6ePwz2X4llCWHVo1/vYRAOvvBCFkIuTqQk4EHpQHfFUfrD9ioXTzr8+4xCB0H
ugxruFvDEGekgZHlaGZisPK7+OFah9JXlDkdcEdDAZpp2n8acquicWNy2X46hhH9oa9SV1rxd7la
ruIUgDA9GLQUt9tZV0AEQgQnMZhAL6sznG1pMGTZcE6EeJwvYzGMGGcQp7zyC0Vv2CQEfx6v8BrD
xHexiETzxu9VHOAzYlBz+BWBRubdPvY2rBQi4elZDP0ENx1EdykClbRPb7fdfrBCvZpCRmH88SrO
xg40FMF4Wxytz9ucLFI0j2Chqa2y5ju1fsJ0IABCsDm1odfaFyfmco6BVuaO8ZWAdDpy9O8gpzwi
qLki7W1Ykxfs5AmohyApe9O/3C+enSmFIg7kLC2KmnT6caEew5rnLaF3rBtpA4EhmrRfdl9zUmDJ
2ZdZZQH6Gb/T9M55gVp/GONBmlfouGZ73qFNAV3HAnPJVnZKhpIoL4AqBcQ4hX/eVVe94co71pr7
2y6hN+0JzxntU8G1ZSuCxDjy5wEndLubWVpMuq7gVlsWHxwtdlIVKqUe0hO4xOapt6PeIhXXrlAW
mIoSQ0CUOHsF+/lOL8hF2aZjJe2gyDweb8FUECafXI52FJ6eHzHRLLIGSRtNs1cNQs69/xtFPfrC
dft3enJ4ItEiOXlvROSUv0f2jSlr4zSO1J9n1/5JY8gjZvCGe/qfe9uvX092v0ArYYzDbS3p0Yum
9CLfeIi+05arINarw7XhcQfa68ujk1bePq6Weamexb870xPyeMGi86A8zBuYJr4wS/69H6r/Ju8Y
0GQ5EWXy9nufH+FqRVHCspykHItMpzcDskzHqVKeS7pU6BYbYlY3lNoslUE7PMBcjkQiwKl5UrQQ
wk9n8RusP/W7lzeS7TD+RI7+iEbri/nYxHsVZf0J0l1mB835PdqtYFARSPC2MLWoAhyhU9T4/fEZ
pUguPeKikpQapOSiXB2xnyNixbWETdpQHzgNy1RUPDDG0aHZ7VI/njl0ddOfd2aCbrJpojtsWQfV
pkpXUhVebEajtKCb54v5qX4/BNMImOt0k/ugEVc+pno1PFtEDwYSlMriFrO5pZpt0yCEmskmOLoL
2HOAycEeRVNvL57BzmtMRklvDe6hnjhsE9UhsrMJWPDVWxvYUXchEU7vmpGj+ehWEstlKz4HkzXA
BfKFFKLWMgS61ImENw3VuA0GdxP4luKbM+5HOx3fNKB5GizMZvwDvImjknnr0Kd1sdFeCAeRdM64
RmvVT9OadoMyRD1F3UKnkfdcxoR8rKuJyqcCBFhj1jVuzlKBLbyCgpkAPaCnZD38JHZ40D2m3pV6
EvVyEktFElodjCUT/iAAVSNR8gNN946lyW+Q+TQiOY640osvHResD6k/4F39psN5obuAASZRgGcl
6GIlQi7v/SDSyr0SGSzqwZmpOlsNf3AbcQv8TPheN3kVuFLYNuF0facSq/r2AN8oLxa3IbCC1j/x
pHrMJIfCD/1ViByY/XEikTfjzFVQxHXkUyNbpctX3TAfG/qSeW7ky9OXX2s42AThYbHAB1mTRsH1
ZWfAQiLnb02u1+oMmZ+XbKMMcixMprt7BkwI8XcR9OoBncfesQNOceUSO/AniJSDF13bZdgLAVJo
r6Xjarjh6Lj7JFLQZ4UbSgrrhU7CLkCrNrh0nK1kNAGTt6qk0CPciRY0L6WW93u4zL3gXobVOdwG
Zkm1XwTWkHUF+tRx+idC0/vU70CaY2BOP7nplq6kRxz+0wtvlKxBOyR+7nyPzybK+lxx+qwXTUXX
a1C7cph/zjDotg2iLOhvamA7RmLIxYElg7PlwOFYoN5iAilcgRKlK90WEUBzB3QQ9/E+pOwsF6eW
UuS9rvipolr8qy0MmbMlpVGVGB2i/3f/T+JuWz7yjnjLXtABkoHCUxtqkWkf7t4QOG2BigAPTRmb
fpRwdpeaTCMs9EVaOBvL6Vig7zr0igl9Z6b5dXIJAE/vdpk9ruhPTTZnEeoH1xOq5pkZcYrX/hkD
UIOvYZifVdYIrc0XohBDeU/uqu2K2h6dCL9fy5+i9TMXWYdxXrAwEBIzqnWqK6uLA8ZQO+/yXDTN
FlVt0Fn8le1e5kDYlTLCt3fE9TriIxc7j5IiJXF55B09RpkiSuCO3MmhTlmcNOEdDP+G2LLqqm6c
wu6MueCoc3b/N/xqTOLlH42No6FmM0PUIcONlbOrCyDSO495l6Mqr5MkYM4sfVP9or1SoURLul5V
/zMdFRKAWfuNOwnqCbQbLMI518EAPRy1H3p34EGG4mkTvgzQjcUIijB25bw+JxwdAqyVTHnGrqYL
Ie1IprWOE2pVw3P/xFP9nXBx9P02kvXL2+sBevZ2dc5p6RFcDzpFaC59g2K2dY6vVM3pwUvPPfG1
nC2R7CDCxvNjRxt6+/SF7JHXCn1SstlDhFiCg12F1GgZ2gEZf/Ex3Q6y+P2Nx9Fr3HFwCkoLAXl1
ba7tYAtxVRMIkJlQ3ymUJwbMYSzmJpHO8PM/7ZViwsjWkJ+R+nL6J6CIELXLxHTkLzI448teA8c4
AMzXueqP8lnYj+ur99cjuZ9N1MlHsJgGmrcQDfHyiAeNN06qSNHSMNSLweB6x5TMpeXKZp/Xf9nS
6SL5QNtuB+CWWwLcqszzw2bP2bVxlyXiDdkvfFw0lJ5DV0Q69IXAnE606xsLaN0NISeqFbrqR8vk
qD2zOH2MC+dGzuTDC5SW6ZAJS8J7aSr2q8Neykl5rQdljVHj/0SOF4GxrK/+0db1O0fvLUjp2IJu
Vky7oCv+ly9tv1pb0ISuXhYf89K1a2QnA1Gm8gLlbEsCyO7raVT064hE4PrGmLBKejj+O0wqDsGw
poko+uREEUzF4wgVnqBlaVpjqjewFHeik7iQmqb/UyXZXnnSc56JjSb2hRdIrSwztkU+e/dLHRp2
iglDdtfd4INP5fWzPazWXWEAMZObOPz9SHXLxZjqR4N/he6t1Paqi37AlzmyK5H0t0QeKSbhJ9oO
4MmdlXpEKmWsyuej1J3mJV1khBaJ8DSTuMzAwCkd884+1RdMu+dP7LSHUwfkUzJ7CRS2fzZuA2Zg
zVQMIM92AF6Q5UsPNljcpaUGVNZ+9wvlG6zIld/jEEeYgWbsSvN808CLcqu2j0yYS0XRQwHexABk
ZB4wTOaJnwYJPQqcIXlcAisHVZDmdXvzwKv3Hjqw1JEdFh9oi2F418xC/0+HgBkXOalf9Im1rZBw
uogh0eT6IGcRRmKACL+MCVMQazC3bhjqOInFk3qFsknebxY3EFwuiiMII3rvQLPinjqYc8taWIVq
hrOMKAZ90QZBg/RgRjbb59sEB2SExPaRpf/tASlwuHpooXzYp1w92Nmh6EyBdo/z7RB/0jhe//Q5
aDvOgdlXjun01LQJch46AtRNx2ZvO0XikpciL/qPWYBnXo7sj0HmyT2qy+mdmL2OrFLCFXTb5cfg
sWjwuWLfdyWlRFC1PTlXdp6Z1O99BXohotRpMCaiXUrRi5ZCspR37zMJjjonCGTd8OQNUT6Rhqev
XiI0o78wRpuLFB2LpdgdWttD77H7ahP1IJSeNAvnbtdOlQZ2EtdqO6vw732wKJ4i4x7Sjb+DPzO/
O8b5v5aBoi2LmRSoEYsiuSdvC60iY/ekqGd2ToAFGPjNULhbJBC7+tfaTSer6/h1Iy5rIZNg2X3t
JuiXLryNJkUXSnLQxgJkiMVR5maDbNTtTij9jEgoEnixMuvJC74q16+rwxci53/d5qVH5EELnwqD
vOcYkF1lfpMAIB6ZILaT87gwPOR4xhaQNh42OIjEnJ4yMscXwP6QBfkebUg9InDjTM3h61NCkavy
pXwaAR1Aw33uDJa2PLhV5w/BdAl1Qaz2RnZo8a4c+/WCcWS/UgeewVJQQhoSzkGpZnfluT0JjOmG
b4jKFZ7AnjIXfv/GLzi4GapsA+RlYBS2RLebWuRqdga1sMjb/Hj+cGRFHb7xo7y737UoDRnauPJz
RIDtQkROF0P1QQcLJ8gO6LhO9AaBhMZAH3BneRtqgyURT61D4sbM/EqkKMEldqb6jykq9RRFT/X9
WmTiNy0vRKNnQx+vtb35WrUOQGVkTod+CbLQYz/vgI1fgX28RD3zeODp27e6o9gvO+iXi/50Ltal
GQHWX2l0RaUg7JkOvSHfU/lTIM1kEDHI7YGsIlDKG11H6x2WKoh9HrsnNVtek+onGqCDbE9PIGIi
RDqMlLV+zbvqvLhNw6dgLSGB0sq1dMOAk4IKnlo8WwyEUPjYEn8o4hujGMwicHw4tPS/H1jEU0Vd
Db1s7rD+YfNeakFRq9NY3cdjj3eDbMlMNJ6i9MJnZJqgYH5QLAmNPaGw/8rJPMRp6ucb7vWxq4rZ
Aa3S3ZvyvzZ1vfR/Dx7zUjJWOzTSm3RD262GDry80uAVey33J0/mcaEZCt8irJNToSULJvBnupCN
R1PtPmo8njG9tGByFogJFQvYsFzjQR8Wj/w8ElNRmlCCz3OMHdQpvo6uylL5bZUK3Xpdvcy3G7Ab
bzSDoBGaBkYtRxLbB4VJjGR398LwtYF4Zd/LakHUrr13OngwSQacLyxMtUJkXv0nS1ArLUn32qHE
1vSFzxZxgOBM21j4bDmiWw4JAQbp+LpP2i53UcL4jEMS9QI+3f0USHm4aAeiL8p1hjpHKBXS0q3G
VcscaLkDK1N5Z26+GewbqHBNQ4E8mtudSm76vb54a3mJtTgZ5jKtroeuuRVOCk9XYEQCLuRlkW2H
RpkiwDxBz/PUY40ZSDRjxY5AusNTUga/1ABMT/BzKuvmp0BeN7+eZTcUx7nRJF5UYO5pAeUBzpcj
K7FbU1IEAmsNx4jXad+5+jQ7Hk1kaJc3SWcn6V/AvrQ+2m7j2PzyafzYCqzGDF5XR5ScqbZQ7c6R
8TqhQpBkaCmyvG6PZ7jsxOv/yc5/gVNbZpQw601GfWC5mzV8tNnC7Zvm2l76IJQBsUq87IM2H/rP
WzxxoR2VMAq7W8+RV7GUXOssLMaWkh58QsWsgwxviKrTZKwW89cgkjuHpC1bz7RbkLERLy5qa4PH
viHy8lRuLgKDuUQuDUb88Nbx1JJsYlteBCzM1ovLJgOtMftoxXFkQyjQy3m4SUyWYYw1LX7JLF2z
mV9u504kuVawrLPp0yCsfCr8epv2hhAyiGY40voGr5YWlE9JiOQACJF1yp7avFqP9MWiu0Yv93dh
27TA40PNpJqKOHrDaNqCtiuBGhCJaMl2qE3SQR3f0EWmsGa8iJfbOBRkLmIyECtZrxjgZ0Dl4w/o
D4dg18xL8EcoM4pv9m4XC6ZYxfeCu64HFGTkq8YnsteK0CZbyWdmea/nBVT6LIoIgvrnr3KZtpM9
/9Dd74BqMREpqFHxD5bp2QW10uJPCsZ5lrFhAEtKIySS0K3LAt+8gbmxElaDW1Oy8HM7tA0vLjxR
XulnMfKAOPJd/6lbRCM4JOx76Y+uB2NswVsFd3e2lUK8c0t+fIhfzYx2GTE+HLo3X+ZNQPIFKUTe
JWGucjjmbfIM3EXuHhtHviKU7OWx4tu8+1kP8lPhobLvf2cNDGtgNZwZS8ERXwkC4CRukXP51MNO
++jh4/sttQBGsnsODA9M4oTQ/zRWb9mwMLQMlkh3O5ApRtS1bMnhpNTSIpOjA7CNWz8xZOhL4oiB
rJB01SyyrstnajlkfURIs1Amw6DvTnzidzz9Cj8v2PW5vW+A/l4RTW0SUa0oJJeN74z76tJueiqN
cNC8T5KpMOgYStGjvHJao27P/H1lgOSsLG0etHBbEpt7Y1frx4zoCaS+MGtK9CtkX0bj+lgw4pFE
JwbwuWkU8YbB0UTJ2qVnviCtGWFZQAUQ+PivtwOeVRoLm5iSqq87CFzZockN1XhUAvwaeaN7gu7W
kuOB62OGCnoJ1GYU4R/ZYnYcDH8Z0onHmP35Xn0HRQflpvO4XFg4ouS/3BGA0NFqPoISRsgCJ3x3
pEY5FwOEhCBGWGV1DJFV2FEbpd0A8QyY9rACixfsYaWtNi/rdPRzDshIndcwVSgoR1IgUa010A1c
FeKqo05Fw2qJHR8VL15ZehQrHIgCKOZtHLCGZMk96BTcqb4lFf/tU5kBAJJI2p5FyseI5zxCBIYm
jBXQRzPk89mWN5cpoZ4U6W1+7Kp4U2abekzwfbR1kvKbGxVW8hZspBuy+7188t5V88LleJ0fsn1s
qlkFIKZkj+wtryMVrf1g2XQCJ2EBL7BqA2g80erDUkP423JaUa0heI0X4LLg7COe/NAGvXY9Txom
OS5R2digs0RAnX/RdbpZ2iG/Z3smF8NNUw3V7eoMEMaLeEiVKZaBcq2KTqEv84bYOMS86JTsac6p
hEBWdJnR57M/anHFJP7LEsTl2wlYiVXe3Efnpz0jfVsC2NFEzgzMZ0pwsnXUwdU4i4CJPqaoHi6B
k3jj6tSB5SflWCR9X+9oJScmGa5SK+PhhfrwRWjoApnBIFYvjzKURv2aTt4ogICiJenwxssXyJzz
zYkirdWqEi0oEeRnO45bkgl23zmCiT85hWPTSIYN5Cta4u7BwQacPVORpJXWkIRltxHTu1/WYF94
carmAkWxnw0hcgLyCgRGx/ywKYYzigIHjCNHEsv8fo9fTXO1xAPkjoxpguPqqnqLXfzSepP8rJMq
n5bq3XGER4xkHFNeKvkkE/OwKiFviasCpVs4uD/vCuIic6rnUSMYjWhSILRkPCuPXVfzgOVaW3ML
mxYo9AD/wC6GqmsAV88Qhel19zgwf6yWYgzzPnJaaMkzV4Dm2CuwVp5u8ND85LV2EnzWjS4MAcMK
jxu77bq48jhhPP2fYSVK7HNtVcOlOb7cm2ELvzCwnl7dcy43FfzqzmICEmUEhY3k2i/Zn4EK9URp
tZJl14TJEokWNA4dzUitaR0OSFYMHlpcZP7lznJ/UstFlBcmdYZWo+Tkxw+RZ2DgN1v9ZyX1Wtrd
7OrHUgRJhaL5UFBtyl+xefb6PPs3FlevOZ4J3tzKclSx1bMpO59+KuxtUCaPEfD8kOyqnxdFi3TR
M6x2cTbYwbYeuzt3eVUjUvDNWcwGZSpCXk0Go+3s4Z1G1Ym5jXrrXZEU5/Chabs4yNOZ/C+L27gt
NvMpduP1KDvawmUVqUtrUfSyR0PURE/QImFC0Q7h/QYruJCUPRVqPtLLhSfdKPdFlC6HCMafOLt2
/xKWbc1nhL46rllvt1JLljH0SH+688G6dNmGXZzTWfufxnsJEIF/Ery87JBCmGN8nfISVjH/Vybm
2B9USFG459UzBusNAJOCGCmEs88gx8Wr9kEDjgB4xD0nIV5qdNHF8L9iK1ZzfZzD/sVFUzYgAV8P
DaIksLQ6GRhG5oEpNCISc4X/0Orm0kFs62SkMX7lwYPRuKENyfsbLhSmO1hpBiRvJSI77Cbvdax1
ybSSRNdUd6JPNHFRLCiP1QL2C6YS4Ko6/I7EIpCqS8nau0zfy7eHHoGKVQTm0Z0DXfmdRYZPYz7Z
b6zCpmAr7nsjpmEuW9KWsxMuLAHh3WOlBalPRhMaLAUFNXK1mRrjovxtST7XEE6tlMpdaGb5mpFA
Egk67TtKxTvPBBJsi5nQA2b4r4OMMNM1FHOfv0hQ5aHcybUeqcx5l7xNN2XrXggkmoLwLDt8FpLR
VxNt8mSPljc8zXkvzXJvtzTNvKfGbXnk6Qkhk0WF/70lsHrkNDY0A9ZLF6erHvQP0VsNKjf/jOm8
VwesJIwWbau6U16OHtAelg9UJhTnMsXsv+vGimyaKCkBC1227dP4ZZfrpihDiPEiuBtCadcT/1pW
kU8ankrNKBfG5GfL860FAwiW6xGyNLEN+LI9DK9mmOOLoDWVGJ8QgkSUrXiRlkywKp9fqgAaIpOi
iq1xdcW1xWStZKH+IhiGiLse91TviTCV3N4JxPTqlMcV5cY74Ee7K9sbCq+91kJTDnZEGC05uMY0
CeKBXeu+126S1ytzM97Im/ov6OJeujJGrbBNQNRuSx9Bo/Wbid51gR7tXTvcT7jyry1VQ/VJaZL7
95YzbvQhVmthLRk6pQbWYcHLmW7Cti+7tuujDHMaN5uGZCAn8BCKSuwoUV+zEntIBIo3iF+HhDr2
HnEeN34nWP9SUjeiMQ0jRLzZw9dikSst2eUjXTBjV+sREQsGJWLLlOa5xEu/BB1vQoNBSnS42od4
JKZNE3aRN0ZNnQeDVIlApYsWRKZ2+IvG43DnFuFT7Rug04//FJl5tK/HwhrP4g6h6/Q5u8ZhnPcB
ec8amrvrU+OC44UyzYUjDtK5C5FudS2ECubgbcpxZjExGHMTRllTXkzKacm0kFR5T4VM2/69s/eS
Hu3xV7jvP891d6DqL6hyGOi1qF6cJ9Hxpupk/wm1Fg5f0pW/T5/cr5TyZAFHcsLZew8wVL9LupfP
l3m6AWKKB1Y425iK7wtPFR8zAV8asOxfcE/nP3Dh6ZI/c8Vyo/ka5fvsarTMLzSi0N1SJDYIhJJ6
oEVZFTX93UcRFWj5P3mO1eYEc81lIMBVyxBka44UCZkQbEjtMEjm0lUHEJE/gsBIrswxactV5eKK
nUwMg0WY4NQufpd6pwVDWIWa2Bv16ID+UbYeTbS1nvrw7OyB2mb4ZhNiAp/g7P7tCq6TM8MwgLu/
X2+4hdg6t2cw4vEQqyEZANT6hH07L98zCnyDQUnmJMpAn9/OvgWX8s7BEK6mkQsciWre2HZ3ZPNy
SxGvKcpRCnPvVIccMMZmcgwy2YmNqBi5Es9hOPml+/c90PIUE6sRk9uXkGbcACHaj2BGeR8f+5xm
L3GYrRJUzIrXHXdnFOGSNL0vztKnpgozKRE2EOdXpJcXw/VZ5MUOpeGaOxS9vzJsDAp4INjt3v0m
UXrW9OCOGtmsz8AFHoHp5F/nkazZUPhftRWn5zZQ9NOxn1wVwVGoPMGL/WibyeqVWZNffgiO4tH4
jO6qyK4d4UAMsOGP7ZzhJwQ69DUuxRFQE82mP9PW6eGJZ4ukynXDZF32GE4XY5I7usglHF3D9OC3
W+joYgIOZM4+cra1PkQMTt28tiZj/4QkIh943GcwsK//YqSrbN3FwA11GhZSW3TqeYZhD/IDztGQ
BQ1+3yxubRNzL/uPC/9cFAtd85y/qI9R8PIhCAC/u+BBzJDapaa1LaEUIitx/1qy4ocxIjty3QwL
Fv3RwnVh2Su/yCItz20CftMlnH5pZwfF9IOb5z4fdc7xrTLe+WORn744sayzX+kNBfcbxnZ5JOWJ
9ETLv4sm4LN5CueF6wwhwn3ZIW7zpzvURXUTs307+GhtBpatXW4YVEMrzxaePKfLdqDVOd2AUEsT
nUlzvo954XLpCgNtC0snG9amEti2SDc6Nf07whyB1VSH3tkNEdt1nT5ceJ491dubRRfpNelFCTAs
8cFK4p39DtT3s7lR2s6PP2f4aZkK4eRKGY9M+HSECXyFbojInm9vKvFj4ss5fAbkoqcWQe9ci2Pa
CFjcEsdz3u7uephyYk1mKdw9vBx2jlnNNzOC9BrcPjtgUpDkdU7QENSMhpoQLeJ65gkuWV9xESAo
2UKW4gJYxrAmCf2+Vqa+DqsEprMtBO+CBD4UwLZ0vn61PbaGQdgxYQyDfhN6co9MjJ+Yuj/PcJjC
QCQs4zlR2dVjkGqBrs89IAHRfnsQVVllMjLstkl6MvBoxyOIaOB/BSW+ZOL3j7iKgw+h1s0gqzSJ
4q75LaZICyOd3NxMlAJK7E9yRfoRzhyEFZ3od5uEOvIEz3yCT4da3bTpyOoFiw/TW60CjAzBCsNq
w9NZ2R5j+X7aBcCqZ+dCBTLpX+8jmOwWCqSG7vh6HmrbYSO6U7mLdC4s9pedfj4dEN74VFJ77f37
F6PAJGyxdK3SKyHp6aYWLAULi/pGT7MFKMOP31MxOLJytIValZ6Wwxo6JmDCcqmba5FcNEevmaJ8
U8laLFuZ7pAk3/5CbkuNgDyEMFirliJIFIPm2NOW6uFaNir4kD44eBYFx8hKXklTQwl6D/lDF5tX
DDHE3+I7NFw27RsASsJ1cc019MM38g0GF24DIRS6bGMagx2PBlGBarOAx0pe3JbYF58n45gM9K9b
m26YlgSsaRrGp7kSAX3T3lIKGKV9tLBQa2uMPoAwV0hWBeVfaFeuMeWtFBmL0mX5PE3+JaD9fQBG
1rAbeSMm7rMKpZgW0teZfAcuOnrD3Blk0oiR39PgR6U4Cgzi1UvcU5oNYzGjEQT7FJ6cNeWVtzPv
QFcxX6FpT15210y0u0GzU+sTPSQemOB+wD56JhVk6tVB9Y6wCI/2h6P0OhoFlrs7iQKhrfejfawJ
NVt/xY5p9Cp4yW5sJBkdb9txXBkOQpGT1lkY3YMfWaBCj68ddyi6d19KjOgBVHfN/YDZ20C1HHPg
7bJ0iofEmJhoY45JjPT+0l4m1DNXrF72Bgs28e0MBw5lJXriHl+HLWJtmobmE4Kwk0O8Tj/BFwDe
G9u0fkm+z7zyvpSpVaRmgbLeUE5t4Q+gzbR5TEsJxU16odPKjeECXXr5OxqPC7ui+8Wa3TrvnSTW
fjxfXZOG+rj6FH443kLU6JAQPsiD11ZZj14u2tEfuycmNs8oubu1DPmZiCKS7UmQQIXAGPPa176d
juqtM/NGZOchv2jAsfKAcH9T1pQXvhwRoWXWHhW0Mjfg1Mpedl7+6qD9SZlrCOTN73t43htZwHXE
nbgDxjOIgRZy9bOxmUZMcRvUsHNRl6eecf/ah7Mct0AYIE7YZMaDg97sZRjDbJZVhVk+msU8V4x3
sVR5K4FV3ziB88LQQ5gAMvWMKVkDYumOKYFoIFCUXmYuuZsI3hexi3kIV2Ld+hGt6wAKrP/55uWM
nYknmuFvW/P5ussVrPEBZrelCpkXAOcRgfU+3+zwn5R8Qtfnb/uimH6Otbc0FpLV4izZvkG5qIGW
nvSxwTQpdZWurv+VMppIFuVa0z8If+xYr1/MskdklsRm0AABvJlpzVfzSiW9wQI8zW8yul3/qgYe
ujiilCwF/8qHI2TePZKNFg5rl0ElJ4WCj0wDRhr4HIVN0UMU+KSVI7BfVpQnZPzYSdNWBmy7dByU
PDy4+V/Lrp0jDltRhrrgdf6NG4f2cUEtvLtU/F4Rey+UYFikCA5lA2V9I7J6rF6uzAkP4i8ka7Zl
FoNLrZGD8mH8Abe3mReuMVm/mNh1PXhXzQQnHmr5FmDUoXNtCzEZJdDrp+WjtEK+CgRl+uUuc7Gm
2/riItZ9qjkUq52zS7VKtqD2KYXfpZfEYY156FE0hHtBxjTSAuX/pwUWT2UN6PuRZ3MCzNTztKaV
KDX03DIYRGIlaEyYjTdHY0mZaUfg4GSogA9bzp/eFssUdQEKvQuLUzhSE8IhPyg/2O83sNjJoaOg
wQ4RLspQJwxs6uygoE4rrB9z8oAe4kdE1DrM5CUhIwMIhkHBuiXyp5yOa7h+Ez5yh2Kr6Vqgk5gC
ChLCXVAT8JqdNLaVlGmokIWMupkmMiiX1A6bAUsOmFCq0HCUMBxwun2jSa4OB20SUkG+H8p9s5Q/
eOkv0S0wkyODLjLF8I6K0PJKu50sg0OzuJW4i1WnoR5EA4OKeJ9GSD1MzLfQB65jI2nNlGDzl6Rw
AAX4zKboEdQ6TrpYcG3jlKgM7yOA1BdWtnjYxBvhBK0rhoxygQkUg0RexgAs1uz0sV9uT1VhCPEE
1aguzfg6bA1IKTXnfV2CvexFzOriCazWTfTu2o/YmMpiIDV2cSkvhEXX/Y10DHC1AsdujjOFs7Yq
DSniY2QsnOuPbMRlwz95UrPlwjspfNT2bpLT+URpM8ohVLL+4mcIljDI65FaKUmW6USmywxgglcq
mjPxVBLE7ULMiTivpnUt3EE/Dqhr0+lsLwST6bhGfdH87lTWBLjqqHxD/NF4QnEcTaEBEb8wr1l0
SwoYrKJVYXLKd3l8cMJ3+nKtS3UfWbaT6cFlEWpk2gCb0V1grbLj4iuwlsK+aLEkyJkTwB2B2MCk
50wqrc4PHjrEPOm1YPFahGzjzXfwsD8gAVHUj8ngqy9Ux0mVJRwqFzoRhcjR9gVQSMxYOZyr7VBJ
/3cEAxdT05ZQld9SatSQgoIRlSB5FmFQCW9DBFrhGYB/6Jy9mDKuY683p/ql1D+ePnPo/ql1OHDC
0a4ovW0hCEfCduzWc8EzsQqrk29t9DLf2jbhn4yTyCNu5awR3sWVn572a+8pur7EUNC0nbha2P6g
F9yoB6o1wT49b0xi+oOqQUiLL2cDPd46NiAqLmo3r4H6pa295NLb+DUbllXmIb/q7WkWeEOhrAKW
K4VC2vOXn+t8Xv2or0fha9V0qoTeCOH2dFAOT0dktAabzL/Q0QE2J+8FxskuNREnzvhL07pzKqum
RO5Or3V2TAF+KiBFnfVBAdnmClF5dkmtfj9aD789dhVg6M691N4L7SUp3fI9Kq9TLnlc/VtHAXBb
9uRK8imSxP0cY6XaInxf8KdKDcRHBcK6FmSvIXrUvtdtl4fC7EMklr+TtNIoGCLgIIJ79ho4Z8+s
q2zfwsaKdQBNZy5J+OhNfxVvxLYiUltOT3mp+EXYg+3tlTS3LZLY+ERTSItTIBLe/gzQeV0HRxRL
CsdbaiztqaDi1EOgCLN6uJYvgXnF1Yj4NLDx6U/cWybLjtg7nMV5R9CGOyabLCq5+rwBiKHIaJm0
RmM1OZifqHN1eP/y0gNNJsQfG7FSlrBC/EWKqXGB3SobPcCqIUHX06Wm9NqTSy8WJ3N8+XV/q4/7
g+qbhvAka+0LXcbDD90/2xabOlloS3+V40ZLRg43SBgmcwqhDPfvdzebRWIzItHMvEA5fGQ0Az+J
wHw4VIiwuehsNIlEay2SecoP+E5nwmpGYQEc+EK5MimDVqy1aKlPoOT0nYy5wzLTNE6skIkROy0b
era1EJdQsYYnPohnkc6RxI0+xg0L/blVKpji0as/FR9MgkTdrAGjpRZgV/zAObfCGWtJSIpXuUML
l0eqHMeAEwX/6OIi4WTN7uhUn09VSCfp2pcuEGwtm5sOMzG24j898hxlMndLvvfauep4Zgf2AzRz
Xua+avkYeQouVPWONhdc8GXhSZVraL8YYT9mZk/3dKoKDiwo6j6Vmpz84ymhaaQrvbbzfbqc7pzb
Jca/DEnd2vqfKRMnyoYiML/Zres6/1lhbCJjxxpoUodgAX4igDB7hFWDptbk/MzzBhCycvFp5eMH
O8r6iDprXsUohddMCo33DhfNxwb8DYBm7mhYlmejBP/dPQRhC4FebW0zJ9XAKFXup5eKm9We7aeb
or2Xp1qZa4HOyy9Zr8oqJq6YRfnWT2h64JytXznHTsPn39HICGPG6QqSvmx8NiA5xNc7r/Iv3Eml
2aVzL+dzlkGEVfi3MiFVUJXWcLkrmRbURV3+p+RG/6AEtrJPbmuQLnr6hzE7jifqPauzaWr/UTfS
vnfb/UOru36JIZ/qepH4rQCVdtsuwrIJ7MC+urX03aI4rxwXElxerY+NzSqpnHcAy7EQJ8ibKsIW
MqnFBJnUeLhBZ5Bw0WgXS5Hj8pSETptTqarNGZot063whYQ1XYgnFDD+rsKn5WrJk5O4NWToA08l
F0jUFLlOdl+SNF2ArQyJRCTeHAAB52cq5/OZfNDPuXgTUjrqLb+Q7rk5s7/l9T8UHjOPxi9cWY0i
0H5pO/nVfSp4lmT6pm8o6TuPuo9pyzh98bNVeSXRehk2qoRErDr1LE/QY8d5C1nQo3dO5McRfu6y
ai0h/cZMU7HsyNyUeLPpjfEBrQ3hzVML77BoPBK9QIYV/aV5Da+mQuoeWBMlUmfZ8wBOVtPJtRic
b46ia5vz6pBpfbtdYem30AD4dTp10MDmqqmQEM9zWc3Bv0QyNNN55Shv80fGX3Bt0Cichhw4inA5
slT5iRtgfSo1JdZunC3TeO7nFYJ0INnfSZZ3XB/Lw+WbVSloIZREJEqOxy52sWwoULD/DUot+Obz
0+OAFgHMB5ZMZypc1ru4zE18t9jXd7FNlS0ZD2crjMqEJ8vXNr7ik/aAkPPHU27ShFsNzOxlfXn2
NYevwGkfvSQ2703usebn67mFXFlZHDz3Q+z/AlXWg+5jNaxAVbNOo/nJtObCFNuWHGSN+EoTzZtq
Nn9/fZN5FRWyegubOtz0kZQxo1t07bZvInYhP+NvnIyXPDMd3YKa0Gf6/0SjZzoEb02SPIrCq0aY
aJSGC/YS74SJYaRaSwEHKYR7QQu1/mPBGlzkCGcXIoSrOs9k97o4/ZMNMY/mO9LM0Ldgi5s8sODv
Gnq5jV+R5EnhT9w1NoNqWoaTL6AppIXTNQu45Un82uqzl88D7AmBzRkm1EPpINgxZHcw2D16go72
lMvsybhBow5HvscZQRhmBFTBsQ84HVWSZk4AkmIvmqPSleO/IsYnqsEy5KLaxvZ0URQq8FRCHN3v
HcoMC/uIgd9L4jmqDBOFxD6dV/jXLgQNsUIN4HOc2kxdcFG9wwELMwjpm/ZKOxMdp8k0IaElrHkK
QtqPRHvH8TDsxr7e9Nnf7L3nFhLVwBevGi7Qqql8dPL9sHmk/W3Jhxxi/t6+QAWXCM2wkhoTcQUb
t7rmf44mTsw0eiFSbh3dbSwcnXUqFQuP1Dp8Tym6VIeXRET1jl+BgLFAHgBB6fjjiIfevCMED7ru
Zf5WAUBWwj8JML6ONdbe6XV+i98gcYsHWPJpQ4GVnR3rJPKtthBBidzAkxByFwZXtqxZxmP7YoOT
ZmleUm7g4gSwJCEdU2h8+c3Bzqdp0lZSbKPyk8Rd6ySwRQTOGuoxJxKEESdXC5KYr1dXjGHZO+tJ
S/cs6HmMRVZCaTkz10HTem4ugvFDs28hTnepkzQ0ovPdJEkxmnJs9EhCCsgGpXI/cnKyPhrn6ztD
O43Px4tdHWw2lmqnqnZRwDdTOVonhyJSYRuC5mSDVDPTtX1uW++EkHcvFEczvJKusuRGxLbwc5g+
CAGDlrMb8xL5DLQpWeYyarY/ENuyQDt7LWvSsGUvJn83pJ25nSkwAUziDalxAyohGPowZm/UzAwU
/qgxUWbMQxxGr34fp3DXISkCU6GgDRnF7p+0gkfEZdMlyjPoKHDJVbgnd8ny6+j+oVgQo1QAQ5aj
CCxp8CVPQ2cfsV7y3Lh2u/q/i7im4/FK1DtKBjDvio6XFyhaFxljlJKXGdkR62KGzN7DbOJHa0vY
1ACl2a9S9K5m+nfVn7vEwhK1FdPrccmkjXe24OxOJ73wfVKzqJ5XvbTaA/3uVPB4qVC+BLv21R5H
2hMLEN6N5heqZrZxcjKgGqStHIxbjXW7PUkIc4xdhXuNKae+MQGJQe66mjG1NtBfBZr+gQjFPQQu
N1oFM2s+6+L+dsHMrRyUlt8kUyILIrfnBuObYjLyMtoUodK/FBmPiVkhtDxIe8VNJJuvhQVQ9wRv
1gvBOGoD6d68QxE3g3KBQ+LTmNe3ui0rj1s9BFgRESfdBikocwrDVtUi0dkuBA8+yftSPtXp8wfe
DlEsNlc0675M+LbalenxdgNHe0ANMQ1r8ZsqCQyS74pIEMm2da2ZHlMyX9tkPkdKDSN332MQR2i7
rZ0phDQ1vZkIpENbq8EGpxuC77zw8q5xzsXpWeAIK2JY7HRPysNbC0vmllcT2xcbINItNjlfEIHH
nW6UNLLIKiIptub+QHlQdBwyFEvO+34pPSULiPSKyDxQ3GButplEXamGEnvoFMOQgkLx1Sd/iaDf
OCvxwI3W9BZLMBUiiVlBrjeAd6X2CIrRYxjJHrM/woRSAqrh5WfBRZRqJPAcV0T7Bp+/e3xprAGk
g9+BlaacIegai7B5OgiyMR7mXqRGgOmTX/jw/Nid0OeTYCwAZDYTSkA6/7aC//6iKPmHDdbVLh1g
108XU/aSfw4oeuXlKXzjThZ5XJjaERevqh9LupH1GGufjTDsPQAPm+7SNIcT6d4/nC1oylVVqAWW
e8XaM2KULMcTJTqceNhe0+lAADZGiIF81nvo9yglJlXQtPryTfu41lNinxrk2/IsjxZq2WjJ+AAK
M5RvH3StrwaXnhN9sFa7SZPaUZT9DlNz/CvdFB2IU5aoYdNxW/q8/jNXT5/KirElyAgq1fOn8bJO
Sx989LbkT/pl22oe2FcchSszKmfatmH86eEm/v9z6ISovO5GRooiD470OvRlsa0nwNLf0sVyZBzc
lWPsT3HexmdKIBxQwXrMhzJXLcKuycO2QCJL4TYMphy3NmPpTblpCkgteuOiAXQ3ZhCrJjScJ7BS
XtZA6Hg/cCr2tMLP4xmE6nCNSCg1fAynCyDhGczMFSmidTZK97FribX66ruVCdGCiryRC7hUpyBB
phQ+ucW5h52o8tcN2It6X3dpMk4Bb/wDY5V00ZApo7ywfxEUOnm6ScR9pDWTiVfTeAjjBUyz9iIb
OCqnZfhu8NfLFbA0MdTYdZN1Vrqy+REi5j23/b53K5eE5AlNAG7FJYCzY51GOJLh0nr87ZWv/cr8
caWFE8qdzta+VC3UMCaEU/Ac1FWj5eW9zCTCX+BEle9kK6GSD3OUVqc3ogthcanb+KW8ZWauBwuG
vnVsElRFNBOUBDuQ5jxeZ+0ae6F8QXgqrPz5ZNohsAWFBHvvatprfPMb3WjaOY2bnC/PzCGDGE5g
cDBH1LpV1orjJPUM6ZXWrpVb8Iv3wS/08UK1flbqOgfKKxvnsgmn5JPxydp0Wr3sflPS62a63dxs
eJp86Zwqv30lo6+D6WU2Eap6AzMI8iV11MGSclSrmMt4rSNNug+XY9wWe7xQf71VxRNlBvZOhe5A
2mkXWWsPLMMIaiR2f+OMtA+qTN3rIkZEcW6g1vHYeLXRSAmGXsM5bJ6ej8IdCmkuwxIqMtWGSqPU
IPTdmD3i0FaM0n5lyIW6K9eEadomiEVupFm/TZ7x+Iv7cbMshkkRpx+9CXdSfYA9nDBcpTNI+7fz
unheVYsXtYWPoMS7xrqQKlg/VAeuOP0Iv/3dOcOqoFN00QdJRnTF/4MuFGn0PGwZXl5pjtFLDj4+
plr/RUssY+ijAte0MGg4udxFAsk2fM7BLwix0ej9FTdHYGgmG7lA6MVy4NJsFV5RpMyS9uLcmgH2
GMQ4PLCLETdNfV1LYVyJFKsy7BmC5zaIEsxjZxR3QeOj3rGCse59pTjaxbsWqeocJbJFEDAhiZWF
D0oE5qE7KVBjGzYHLnCARchlErmHOUJbWL3O15nUeEoitWX+Q33MN8/+PY7Afei+o5MNQrM6jJXx
gbooOdU3jyLWKtsCn//vdO44iuQPnHY70i0scelL0kAvb1SFi7fDT3MY+X0gdfMn8W5qmQSn05yl
GjLaouHeB6c4uYFIc2pBrSnOfjusqIJc/wEJlX65OpiO4/j1QTmnaRRfI7ITqXsz4O7gRh0UX07v
n77Y9s5NHbZK3bmUQfwkJp9auB17sCo8f0EJl00G+A+HvDRMmUwB7VWfcGiq94sXY2uSLgjOe8bu
yywbwDlEZSyDdqQAK5HaJOkH2u050BoMREi3QY6dp9GK+gGPGx93CArTOQsb+dy0n+D7VL/oWZN9
QgMxz7Rs5q7HbBGyURyRjaUATu0En47WZUO5MKhRSeAlpGl1wDIykYN10gX3zwjrMjzybFYk0uWB
BG1nUWZiGwVCg3WBTL+pAb1pB5cPhpbqj9AccGcZPm8XjcTMv74/RFt3p9ICcJ+ws2IPTe6GdCef
jY4ZZEJ/uKmFoTivgTzrM3pd+9eQzVSf/DTqtCsDo+GpjogUjxVrPe9hGO47vrKoYmsKissJlpzt
A9ogRT9uifpDHXRMVkYIVTD/YeGyHTgN6I8Jwtc+PeMRhUxoiD5L9GwrmCU4LbQEE71Ji4zUAtEK
5AkQmCYewQKOwmSfykJehZSP3VY29gRqHJVWdG783fe/yebe3UbYf8iZAXx664wunXj9igwpDlkT
DSyRjGbOoAM3kPpbwWziceGbGvAynYKOR3rufA3hQoUdAz5s2x5kPU200I9s9LoCYsm3++tU9rqT
JOP6k+gC5gTO6H04caSih/vBkTOFnI0YLO28dKBeJQNDuYOCCkLE2QDIdiwUgDnnNIWVC0+POzHD
hFWbQ/ht0pcSda/osmfwa9483Ako/VaWCeGfQHRqUDE3qjvmnSsWfd6lCfEGdD+yIkBiho1+b0c+
y+9zUpu4Lp1TLJKXA4DX+wQxYyN3pWpW/TGcrashnZVMhHcUSWK70Qr5W5n3gnfhhnC9fmPgHHP+
lne3a8lH950PC4VDBJ/sRB/ErjzcylRNGHLiV97ZPKGnCORAI50jNksR43vcNVpvqLfJNNyoOg/Z
z/iF6K/ZcOSrIXa1SSk3tk7BPQRnnIg/ETbbbzwd1wb8US2nsXckGmj0tIp14QwdjYGvAMvZzvE1
/7NIms/jeZZG5bmdpXkKVk42Vf6tYx4trgBai3gs/8dY498dEMF+NzLE/QubxfHNy07DjnZ8/DGd
XfsbyF7iWjNJbZtNKeqYg7i6vYHuwvm4lU4z8bedpdrj2gLjWXnikQ2LvCuoJ2l9OtjDDXiJGuf6
8j7Py+WOZN4D0eC+FqdulRrlhasj5ZW+xNMcOt/esIgo6feKX3gEG/Z2jUVPP2i0HZZGnOilUb33
7Xkn5m7pt+n8Ibu09zNbQv6aXIqAKo5ew8ZjBKuUCJ7lcbV3JD3oB0uynTFH5/0laqVJFQAqd/Hz
OvUDwJUPv7K/ufhlNiL3x/IuHwrcp8DYc3ygfdYPdUbUgpnQQkGm/gfZrsGwcHjgfnMZCBa1p3pA
WzSBiZhD0BQc4gGxqxFGWa/XkzhPBYMDNnp+XBdJ9Wm6PiQXlrH17TlVsgQ9z3CDYouuRUsuyO2l
sY1Z4oIKYs/Olzbfkh/OXcf9ht9jTAyy2PdJlin+q3qFlydZRuN/6i9Z54uLnoO2HqJOhRra1dYD
DXotN+jlofuZ9QhWAVNpZD4bNne0A35RsdX3soYfl9YSiOtxuLYgS4JhdghT47x6F2MNEO4NmEwu
C5pkQVUMyxkb43Zj1I6LIFehP0Ee1Dp308IAmcC+SgUql77Ms0lV/ZD/pwy6zkrxoGsvdGO1sMGp
aSFAQcsF96/B940O7TbyR+pj7pRhEFrBfAGPS2NSOdxI8hkZUrVakxY6IiMioL0q5Bz69hdsktvo
SJFbF72jfCzwOto9UcfbO1j3eI/73tnERHkCyYLLDoUso6BmXy/pi0rEf2LrL7+TQ4744ymsDJYH
H5AqXHNBoNVI22XaKWLBDm2Vb89799oSvU17u0pY5YS8tryR/9+vW5etW/BaP4RAZFsMp6lLrvzh
T8FOaeY6lJpOxbT8BYNgC/Wkkqymn76dP6bPYlts9D1PdIXgrVsw8XptIA8hknLDtHBxmqjv+92Z
+vig7cTl6mP5DOrwiCngZUjfA9Z1ya6eOosfE8ZtJBw0j8cTGnOMDuLbzYvjHBE8Cy7LQRGzJlbj
+kLfLfahg/o9PgbgeVtnxISpB8qTcom5zOWJubRJV3g46gq0m0Ky7WjIdGo0iomG37MIekmANVOY
uC7eTq5Dvzd3R+65LbJKUxlxEMay3ldoB7xW2vjKiVt70mxciZ+SAwsnouwVJ3OpEukx9OrQ2sGs
JMqsjtFxd5LW1BY3wyYlu3XDxmRIMyBonlCRYnhWZlUaev7cejrKRcyEswDQSo2BrXz+weDTwZj4
MhQjenyj0YPF+xW2Xlcs0q5M0DwsrOnF79KgUFvyE9acXiPIHnMpLd2zmw7oxK+265c/H9vgE4MT
qQYs7+DwxxaBED5Lp5uj3qz827paq9Qem32aFvkqUbQk7QieUln13myAdPOQGPjH2v4Nlt4YviGj
r3VPTaiEt2xG/LWrJXGW/PdSUMUwOmQGQrG3HTb0nhaCx5n5yXcN0+Rg7/jYsxWSTB3M6FW3qfQz
BNEAI/krvcG+Yye4DMi/pQ0XWvbuEbPx9ofewimQV0cBRVCkAjAEYTwfD98xBRj6iyHB09M2hhSZ
/ohke2xXVVqmNPji2cBk9BiaRqq9G8UMGfXUrRjgEyWbcZUlWTE+nLqyvjVu0poc/vceJNj7ErHI
wpvxO8l32BHdiFecvs4v3yggAn7FxR4ypZqASTw2/JDPn4+IkP30y7pPHFMSfprLYSv1GUTU37Gu
Eaaikgn2nX3idqSZU+v5lX9f9YXtEsOI3NzvdO0k7zaHZ5lPSFJAjXJrFbWoOxYVvYwomPMgq6DN
r9cFhsRAbPm6/WxxcEX29Z4ADNzLLJBdqCyWXu9LDiGDtFBVs+JRcFYJ302pB684ENMdfE4jHhqW
/v/yKZ+Z2kXvSzCCIxTJZxO6mVhvKxcQfcB0MkjEdUZJ/GBEuTQgMGZLZ3JLWSA0BZDJupNIfMAP
BuxYBTQNOABBv3c/XiihUXkTLfof83UcHCUwwKtZ7JcvAWgAjUQh5welnO5lkXRrycLTFWvIwZyZ
WrU2n5KEqC7Ukc54eu8vnYZ7yYF05nBxt/eDLPpR5PswOeqLr4P00FyZnX7bE4w1lxSAp+1CWwV6
Je69rTyHiG/O88s4gEHk6NCl9KwjnkZBlphblptOIkbZkoCkpe9Uq6x06/hKVX6U5NGGGE0r/9IH
DjKCfYAtrX11wq5Y0voKmBo6ixQEWCwcLuYuiP60X9v3EGOtK0zMwoF2wY27xKRP3ZqL0e98EjJS
PaFrq8Ki3LCGXrHCdGt6EGbZMd2Ag7t5J0FKr0VO7F6b1+0nV1TCz9lH+1OL3QqWHCk5QkRtFurV
VP6Z6UpFz9OOHbWMsFq3gRgatdAIJcjijPj2vZruBHkIgt5xaHOVf47y9SJAXVm8+HkN9Cf9rIR0
ymFo99DOxbq19TdI7gDOWVaa6MCVVIG9Vn99BeRj4pj+NgZwI4HOz4xhloyKV4ka9AJ9PPrH2cFR
oIY6PF31d2ljPJwgjt20OKBZdRada5M2MFwVzzK28Y5VJLzsHScrRrAcuEMxFVj5i4tuS90o+1io
UPlm45oDZ011xYj8HCSFoufDZE4oJCrX8jqyY/xlsdC1hEtAGbcAuWQdIWYWZc/NxezLjrYDXEO5
XcQU/L0C1fIqrmx71IbYzHYbpDZmbeDFbUffwzV4kmXgXqvFc9hUQVYbYCaTS06eP1MC0beYoBjo
2ylcb8Wbm7/Z14FYTWLyuRIT59wCq/x/iGa9RG+cDAEl50kJIY4WpGI4fSTpTToHJgznzNGdN+Sp
GYBS8q/LHrONzBScR8x+PgP6autrjklLYMso19VCvjB7TZCG2a25UjwNxd+TJQRZzX4Q+ogEeCT4
kS2wRmb9kvNB7AlZsa+wkQfkzBgYJni5n5hbD1x70LaBJpMIdu1XloLVcr4ByQZYjky/se5Gyvi0
/xMvCLw1AR2TUVLXU34Iz6ETAi82TTp7zRuLNG+xHSxdgy6NoiivX2mcrC9aM8g1iRYZEPIxesUe
o52D+F1jWpnb5s3sijj9zBbZPQJwyA/+TZLwiQXlVzG3cLQ83CfMfeqhtX0Gw4lutA7EtUviTSbX
VX5FnFZ0q3/O4vhFKeslKP/6bl3XVRb9MtjpmYDOYNDKDUI8I6qdr4zPPJOoSpHNv9nPb21i4IzD
1jIiVrsrXJ481E3W64CeNdwrrDNIK9mqcA7ILeT3iSYhKwMoDW4zBJkH5ugXIP2Tu9PYPrKedNT5
W9uUG7tlBU3ApLvvP3SVqfiKVIulhxlaP14n0IS3mhRZWTY25HQOC+HVT5WuP5qe5lzn9wObTo/o
ZanLlNIryAZnZWaXeuqj85Btw+BriqMiJCIJAJBgn1N4+YbEXWPEgoN4Hz685WHzJ3p4dU0Vmok0
kL9ntGWPyXA2rznbjTqpSPDlODfGv+0YncBaHCKcuwRS99+df9e4jsqBypI5K7YlyXM+HrCdqpG6
huCnccRGSPKo4lCmWla3x50Eq2sPJkNqgwRozU1gAHZzRAl10st0iM8EqyJRBCf9k2jKY8INHbm6
L9tIZHfvMCqu1wPKqPjHUzeH/rBtAAYk4475RKUacrRkBytk2Zj0nbnP8PU4+mPPtp/IpJk+ekHd
WXnxxsJEw2WGCt9UMuKl3qP19t1H/j35w5TZmkl+k6yfs/zaXlcNMh+B4uvNthbew/T/f244yz3o
swNZNw0swTx2DanJ20guaTntSqsbZMMOsSeguxJr7lkjOplJC6hldjTHDunCDZYhbtFXClxaNo3X
NZs5ceylf9ng9IaN8CKNGKyAwFszEy0+TN23A/66WnB5TfRxDFQBIP9WJoWwX8v0QbevwRzZsw+Q
wlPbEbYC1fsVsCb4lgmRzmLZbn2ymysCQ0V56VjtO0UNyQ5iiEjeRL56KEubI7JLWk6HUO++9Nd0
Nj4QZtx/mXgYY05brDtBN1UED6efyGLBpcIMqpLR978WwUb3LgWzsVzZIiwQ3la9nSSiEEF4FOFK
3ppZnRVQ2YCQcCiDCKnoQ0FEech38JdGTOugDFS9k/2I4Q0PbVaU2bcKB66Tj2c2fpcuwIWvTgbn
mp8+4KReCARADPOqW+dsElg8S3+HBhxaiyrCXZAkSCI6sxqn1BEJ+xSNjlQ6jZHhjqzlpGAa5dPA
QRn7+MN6hhXGTEgjrsrLlegkdkRoWaRjRQlF/4nn+vPx5Z7XAHhhiM9ylVb5u/txbPNTIJ3tlFHa
ruNC7DVXfCkxcCT/PT1rtal/UwhRWiMhc05Ly175ahC/ropKSQtoT5KcK2h/6XjH7xEtcBcw6YYs
1K+P+IVbol5eDbG1dD8Ti1VmeZOJclZXxl9kp6DP4gcanAuIO0uUmQyT7JlyInUqbsZqu8huXzEn
mEeGhZGpHsj40NKB0XPBd7DZG4ZfF2H859Xx1YySIkOj64d/fIodGe32rYVhP/Hi5nbEOKgPYUe5
lbYXKjdFil/Ia3hOmPc/xolPCxVeXl6z2fi0eDOroQNDEuwcAH4A7WckJzF3chLCMFUlDDuiK1sz
Oz3eTZtDJMVs/5sC02eN+x4eBz8BKBCysyExIyLN1BaZWExaxOpmQ79gIz3HuJvENhMe5/FMN0d0
isB1jLJ/U4CK1wplCfDPQI7jP+T/oDhhcEOmwvvp+KODFqXbASemhONhOUaVgJtdoTxkpLhni10T
SUlDr/esTJG0w44mF/GBwgCuXci3LF4fJqaOUjKZCQpVtnEUx0kVFZ5L9lcr9A7dzd7NhnM0G8Ek
JjHKosqo+YjASUZFnLJNjErTt97v2iUi/wSIs520e0rTeKFpgmHkSDrZhjhxJ45OGZOag6hU1sZ9
xOMWopzkPTRgprw47umhYINmcr4Lh1aQsV78EgtB0rgEK1x0PTj62gv1eGxgqWORl4TcYtXDAi6z
cnSmuzqpDocST4g9kJqH54NzykfwEA84UOAWYlqnQhDGnjGGolkNouid2nrqk6LHcE4bINWE7EuA
KhLjUTcnrJct/OAR+fime79kqGN2XUtzRaJbsC1p+oJ6PaTY/RuaCmmHbWdNAbnKHKPBiKymwslJ
cIppQhj6V82FQ9uqVrnS43ZpwBNepZr87oJOHEPQvXewYvOPLsikGXDpFHqgrnHk7kZ85VMGkok1
HyF569ldFoo4VyCrOV8xfCeG21rJK15Kb0WBkR+AkOlTYfSPF/SiAXQyE9KTUFSCSwKm/7eKV6R2
at2SCCKJgwnIEOhsrRyTLDlGMVtlYbSdKBw7U8R/C5Uadu3QASx1WWmRHnq7+eibmzsCLl4nhWFj
l3wxU7wl+gPw1o2D+B6p7klT5WaHtVblQxD/5xH/zoqk04axe2BBIfk90+eAjL0Rw5xfzBUK8h1x
3H4fy/VoyQ+KnbW3ZjjZ2stmSvzP7kYbDUgXVfU5NOHNHGDpS85YgQHMBopSMo/gcabRnRVKoEFV
1DNKAiIqY9yrAQQbqPMuA5YGFux/1eGeQjs4gjGza9HFeeZSlwRdrvSGqbneCDw5xz3hHkk9ta0O
SolYWg0Lpi6o/x8pYjIIvKYRRSsIT0PG0U78hLTsvQLUxF5gpkDzdEmxV62VvcVV0dEIf4nzC1nj
Ac7xUZMjLm7j6NKYuOB4CY2NfMujbsUwFq5+AaTYIpfzE+fUoPrk0ZTxP1NEoubo1ZFhEUphRsXU
ujjIMXXmrbE6doZAyooNsHxvfgBT4mIy9KRiWxua8humuQbT7Z9snOcnYl9qmu8C9vcmC3Z9wP/U
jZYX9VB1abIq3bUqBDLlIuCP0PvRU1QxR5nS6bQR1Tbj1CtPc5cf2nVYpZCaWkpRBTMq3kN0OiIL
FRJXiFS0JVv2H0jZDYnarcwfTVVIl5BXV/ZcTpyXIAXko7G28y+2My2H90cRzAMXyeUkuEh4K4yA
QTyO4E4RCJKHMUMQOTErGDEIBRgsVC+kZeSNuhzvgzt7ZE/k5SkMYHRWizOmk0d2bkMnGARsfWrv
yVbe8MsoybdIFaaGRo9Xq6ajVi3TEmgnNUzz4IY1TtnAq3YBxN30DH/e1fkCq2/puCPU+jj2HKeY
3ibwHC6xE7ibvk0PLNaYuQpPem/Wk7YOs3am18MMsbsDxBnpfhJdQA/i9rbh5lwYEo59uSN2cXpL
ASmA6N5JblUOWOHsHvZl082fivPiFP+OpjY+gB6yRAiIkCAXNjIeq5T2lULgqpd9EWS5o3l4KL60
9Nx8G8V8ymoc9TDn2ZXwKRLZYaukDtGfaj79TlV3tll2G0iFRzrNVkRngTOV6xtpZVxtmu6uXnY2
Ky5REsIUEeKNY9MNWza/6NDnzxK+rUM4mHBBP4xb6xkuKuYwF8qJ3Z1+hzLXxCDcAkJdZZlpvIgO
L/DmxnkDrlaOEvxLrXJYxd7Nxd2O38q8Y8yTSaf5uxVrda+fJdmQ4KUaQ5YvUh8OOROXg8drT9eK
myGI6LmcfUlY0GvFv3TILuODo9Y/2zhZIRM7jgDRRCL5FaK5QaPRw12ruBl+XYkTka58ZfVQoOmu
o47WjONEUFNdgwannn0DMAwucwJCIpjXrv7otQInXWfLlegArV9i32FYuvpqc1lX9u53/ev4bQ87
heRJHjhmRLo3CyuoAgRnSuw10KR9Sa5ehYIt/aEuXWIbVna2mdl2QaSACBUZMkp1SuFtK3asNcO9
kTJwfcnzVVFQN4Llkbt4tu8K1Fi2UZZGxg3s9Wcn5VcjINjkboSE3MJCLGkAV64jL/IPXUozin1m
yr+L7vBRm9Z1HC8yrR86L4GwkTYul/Vgr20dM9zAUMWNqqufuXuQ/UhtwjiENo4/XXzLpC7n0KhW
vvEDFNi9G0w6l9svrczrDJNatxXJAT38enUqzMkZFXIsLdYbYk3APQLANt8shomfGfvwx9crSQGa
MT7jmAdHAsrLxMAyaBF/aJ4BQ4Hs77jiQb9hYMuzB8n0+NjgQfFZLhOrEbYiDIZLmeMTiAfkCk5r
+UOEIhYZaYn7FsWxJ/41vKUCj6cp6iy5jOPGyFXI3jWIMJFv212YcZ5kRiPwis6IKQult+jWBQF/
j6w1MNfv2F5X+qqc6FYCaLhVcEf7PRI3CE1xkvmFg3YWonUAYteHOcLxwVOYWFopmDPd/2P9TI4d
82qGvvn+hJQvt2J+bAq+yf+546N08BcisAYRqa4ylA9KlyvJ81POc+KFEZD7QW7Oml7OWu9TCTaJ
WoO7h056zDjXB/FEFl2JFHuU1mvZEJxoe7Uy6yC1a954JGsqy8wvN+jjhUUE6dM0Nr/FRAL4dj4w
Rq24ukGwVXlyALGvj372E6AHAq1B6MZoyWRepwiFDvkGic3xkgfgTIA3EnzGx6hhDDvbQfUXZPw9
7GPmeeG4n6w4rUv6a8pUMnZ0TaYBmlXhjt4HA+ZuDHcLzM/akiAt83VnKVQCZQvi+up7j7quQ8Vw
RLBCf4YymLqDA25hcDYW537O118OU5oT7TSTEU1OGEjHyduKTfKmjGjN4m1icsmesBPLxIrhUUB8
2mmquo1xn4ycEuDPCOYQcx54N25z5o3lZwvKWn2LsDO9/zgwrfY95T26rmQhQW3g+nsjQs37DgXM
xpzB+IxveH+q8gm6MMV+DvGf3eWsaD4Zwl4nKvBAwrtsGzaKLT6f85G1+k5vOmJrfHqGhNd15aLh
WmEJol1X5kL9saTLMypmuqTe19QGIrfjP77Jcv1ukrhBvzJMdlSH1OfEReGXkk92JLwhT9vMS15N
VIQWpIoCj37MEb2No1GBtCy8gzRrvo+hg94EuLHETE9WLFsPslbkJ5BkvQERJQdB39Me9Nvdm85L
QlKgNHty//WAWWMoUNjbTaX9ZpdZdvpQhXk2t8gzegOBCEm1bA8c0XG4O/rWnCIhICo2UqLHeex8
QX2joLOccj2PKIT55HgnjSyd/E2v8RJvwRn5T/MshOElTFH6EivsA2GMRTk/c8GznrHy1WKbSpZ3
JK0x1KDizFPOHI6w/7UqqKt2Z42pqfMNjh7DbF0DYh/mEbQZ/MiAee3eqh/JpgouN7ye9vMZGotJ
4miD7gQp+wISGI8ylQuMN/CrgbWr5CLIoWpsGbH5xu75HpKVeY/dfdvtxngNOrUwCYUdZc3l64QA
nD89O9rYAUOeqitTR5XtQAI39t1JQX6aIctkdTesel/3z3NEOTKFfu3RO8aW5F9QqebxEZ6aH0I0
uVderv5uvMk3mVXcdaEzN5YxCa+lFnrQcD3Ul2vg0PkIDwmLADHPhydeUuzgqOs2m8JCVklqfZ1U
DpSvu4r3lhq6xZ/Ytv6TbTSW1nOwOoNyP+GRpbgzjs/RPGxaYxcHK7i/odOStxboitLAlT/fODPJ
kbvaLRD0YxtcGuDEecFMU/q8uK+ezMcZxvtMxYtWpr0GVHVpEGVWjDYgkQgmM+c+BXWmc8wJczp3
8vulS7QM7/rslKt4s/kPRMzaeNeyI4bPbfHAbzUWgOZGit9PV53vwQ7o2z2Rn1qsbUeVEsQL7GN3
OyHBsafq0j6PLxU4rPpX9syoV4tT5plT1ZO6QK2dcLqF+e85O0h591NsCPaXSY2jhgCPZfrCqslQ
IV8BCXlZsY671hl1ZU1gXTgNlq8/WV4h9CqdvwS+lCAXi29jE5GOCxFzAcuxeUMFJwkB+8YhqXdf
cejz9kJrVzcUBIJ7Y+odIRul9vCTS9SzrjM2d0AE34JIykCt1Fr5XaTRv/kXKIZDFGuqlS8D5rAp
ZzHPD7TSjZGrG56hYxUPl8Oywdw48BS1KncP5Vf909wSPblMviD1GWktBDKHspkHHGMoltGind7A
je21KCv6UXZ0a3QR+DA0T4xuLCiM+tgQwvc/1n7dlGyaHcHfW1OgAEIF/8llHOqqE9C8sfZ7UC6s
deBVT8Fnn12R1GMi23BQzGqTVCbudMnImyi0o8OqgTnodp4EBCYaTxf+w1hDdqF8b2KG0GUU9O+g
CGrPX8lW/+9/Fw+1T3mKH3LBWEq7jAqPim7cZlMhUj+Yw7uNr9T7PCD/UBNggzfSka6yhmKnMmyT
bWXfTr1GqXeQJjFvdzCUKCYMaYltn0c005lmLqlBj5J/a1hq+9Y3COClMgI/Fk7ep+ucTXu+zW48
5qbH03lXuje6soABY89SkV+nsnHHEmDnCUNcLTcJcJTJMYL8M1ZcUxjbwAhdtY83KVZdkuqNcViz
gAow9ivfZiz+ty34utHKcB70V13TRXD1fvYzCvhg9WW8odrWETWHj9bSLqwZAiI3+3asIznq2ECL
vx2ORQehpemBMEJlruiY55fq7aNhCOqg0b0oxnAaZFCxh8bRJjmBOoGLBuPcOi8cBJYKxUCQi6CT
lHF+j2xoQ1AcNr6U1DI4Fyj2afK7az19j0MgFHyuKxkDuzhCt+PapGrkEX5i8V6EIPXLIiqZl0w+
A9Hkd19/BY38Ys1k92NmPxL1az4RuXzPPZTrCPExzJSbX3w/VmX76HgmMb8ExPZDMfBiC3jErWQG
9LV25i6HEqzYJHxnA+YDx5v5nwVFqcBqPwsyL2jsQXTlow3JsT8mpeAyK4Ql2YR8nOKeeMHxTfIe
2tjBqkhOCWDnhZ6w6YRNriuOsz5CfqWRvgxQ0R+gErXdLl15Mo29Qltyvag7JsV2SUbwf9MdgHIB
ZfguzckxLRVawpqUKZhJeYHHMDxSH344qJmIx9oe1hgMVhZDvFu3Nh2nxzu2xgAcbD5EYxAHtTjD
RL8rkQ7txD21PE4tONDX/0Aikjk1H0nlHtDoysbnk91sY0XX6BpNGHt7+gkJ8e//2mjFxks1ILcU
81mpgx6mvXsZ+8WN/Rl0LBV9BNzsx2FreZocBffTqJllBCz3LHnfGQZdcLBYqcMkF/RMBm0VFbMj
0rcKNYhzfRDLR3omYcKzBI8K/k3xcJ5+UaujmrkpVhZU05Zzt0NpUM5KNjURcKOa3EHbSE09zkiU
ymc5nNn6oAxYvJJWJSQ4DkhRi2ugQum8i40obvnw/YLqzuRlgxGH2lFajygtQQfwcMn96cIHt1vW
8k3031FM3nYKx1Q22K0DqUW/oLR/rmsqf1ficu4p4zLH6PIijZNvel8EhcOpcFmUkIcez8n3Q1Zx
K7JFFG/pBtfPAdqQxpMnz1Ajh2qBEaGBAIefV2X0d94vLN2RYSNIO4LTiY+v5vowPtTdWmH1oLLA
XJsBkr2BaoMBvHpiVLBdrjcEkzbjEowFsxURgJAe7rPZtSDL2xt81Zb1bE+x5wFxg+oPnyJnR/dR
iHQgIyc91Iu0OuFP0OWaqwOSYgIQHLhr53f4lbrDjAwJgqO5dc0VyqefILfiHYNPVtJLcDfUtlfT
sVHW1uPqagLN7ER1Rjlc67wrelniufsXYawOIWagUukyCrD0ckSfQs1amIxd99ZTKhB4gFCfz0Hy
7tkWyRAxP3kzrCwBbmazEVllpExXzgKcGafLJ1spLGeiXSHRU/pPFptaTBmcdblT6IIBxB8thJ3o
qoRQbjBSLn6MH10N227zc9ZkHAQHd5jKTz65OVBpNr6kUz/H09QVVh9hqVxj91fnGCSKKlDOgqnv
UgYBK0Fs5ovskaAF9gZQr7w0ZO/t3EOcArtUQWMuxe0ImE9quQfVo2irLHCBTH9R9ZOZ0+WIENrW
n6VFTgQc1T/pKgeGqjLPhVpZB1VraehY6GkMhOuVEtqmutJEfnzgUm1Zg+sGRd2b9gjkPOLXSrxA
lGt9NekO7FfnsDbD2owiaVDpitzjkYwEMbZfLmbxKIXWhqrpF3NvDie7Z2eMXtjih7I9uapkhjSA
y1DP+c6Z/SBTXFTb8+2AtFKp4+s8Ut6MXywSG408kMxHqFOwqUUripZuJkAm4bp/C4alxxFEe7Qo
JMSW+Stbwx5TKlTZdXQJnTPvGqtvnLrK6AUGONmgV4Cw01JfL0SMioRTTkt+RTANDxaz0Zb1vgvX
aDccD1omC/tkWzZqjhks0CT/iTuogfpt8zucJKUqovG4VSQvrnMd80oDFlMIFPaNKj/u4wOWZtp1
WoFHPilun6ISWHoAY3f8f5I7v5nbNGs6Tubwsmw+fsTQi/INwzEU1jIYnnrDOf26asdO7i/TRTMH
HC66Oox+9uczziJYA7oWLXtlQczIQvMhWZbVIXT6qK7XkwB6p3WBmVX2dDcVg7TGX7MEblTbJyLx
tNmQj78dj377h3BBR4IQI4zhDNrbJj7Px3ThuPkFJrwU/AiSmNHumZ4LFV0svcV0T6oakhz2OPQt
1fpgSR1oPjbBUCeh8d/oQ+Aq4fLIcu9h8aKRPt2IBcw9P7NosMi1jbmfmRRW31sE30oc64QvWoxH
uATxDC3UXuX0z6Hgniig62lIMjP80ydV+YQMkdY0YA3h3YAIyAcJ3ftzwVN43T4PS+2EB6i5Yztj
X12/lNxOOYvOsJiChrnY/Z0lDyw+JVP3CI9nbyBf+/gRb/PtONyiKxORDBu2I0aMyckW1F1qT4jS
r7upxtgH2yA4qsqhldKhwwzvFR9GcXCbLaMbF117jbgCyRq/btwF4LEYDwJsz6pWToJZaxrn+hWu
ngznCuOylIkWLMAwVwqTsF7ZgrWTBRhBWKqCed0GJyyF1yJ/nEC6dHBqCqEY5C0JK6ex+CbNB8jp
I9dRE8qfPBro7Ry57N1GEOLmkDQUoy3Bka1p9gwGIKg1BKfRbKjzQWxbNkxdqhoVYLeP1rZCTxZr
EcvjEohx44ENGnvJUQqNe6xu2grJDZ+5UwtZ2SxNFQ9CTFJj9iU2eilQiptClefvJaFwhLEahcAc
x4aQ4kcRSURfbGIbmljiwruReNSMJivRQECY6Rl/+xoiM/tf3MGywtq32qKGbxQrnU7+OSfw2SSG
vTNtfe/25PnlciR0Wi3RwErgzUeTqCg0f69uVEKXzQzseBgd97O269p8l4WSaxHRp8EFtHl9MNXI
adqyGjm77mPMCxlUbEpkClhvbFaucBZLHbnEzTmswqomBFZT/Edz+F1Cm/iazv9hh69hdqN4nmsU
aB7vmGrQaUTMeipgEruqIFYSDwqT92kS4jzwMTRMZbOt7IizcECeRY+ROn0L25eQyfxaAML40gQV
JLWWGLcezsMJy86jl9Ue3z7szGhbmt0oPBsTpDe0GP4WSQ0j6NEMlduqCj3yM7URP5zapwaYXvba
MASEDVxMQW2L6mWqsbVQzKN+4Y6F7Vu09SbFp2gs+pcEsUTiibdrIqt5uKpl8shfGYd+7ka+OBPj
EeHn+5clAP12STK8/4PQ15DntZPCl+1tIVss3SMF+m637P0InmxubixFjKSDjbR2o0DU6eO1l2oP
c2K5Vl5H8jj6mjtC8ZyNDhACE5RzLPWMviqNc+URQZx3RDMZNUTEp6JZTWKeUXjhTcZBBivc+J/Z
FgisRz4/kWoDAVXsFqg7CjjXYQzdCXfWftKkHnJc6fNKEzKGdhE7UDsvc+NlirqrCU62AXCQx1xB
X6/8u5TYUPAVOOJ8aZzVXzJHvDzW67agV4E5sILsyB/yDz0mQLALQ566GZWOn5oC0y0sn1qRvHGP
yQBaQIeEgYAEaZ3zPTBdtFgdnWu9Fqc0oumlK7GesU2jx4/SPy7i69M14cp52dp9LLfeQH9iel7t
aCIiXf2H+J29PfT8ydZvNKd2/gadu7J2gG37Ir58/Ouqw1YGXmQpH6G4Ovindq00Eh3dHJIvrkc9
VpB1+DvH/UfaIM9KLo+HwmTYAtp6r/kPNyupl5FsVyDiimNEPtuqw3D6lcMkPQQQNj2eKIo+AUK0
dKpkscVjLkqTplhyBU0NbUuJaWAI9WGIC121l88F1HJ93hQFMVXapzHJLaRZgMqsrtABI/OTKdTM
K1MzrdiOSEHiIq72na7pBx3QJxX1RhUVKJzR5+TsTeTwj30dK4hxXzzt4Qm9yDfvAJ5QChHj+1Lf
gnNFE3c0fn6ubXSpjRARsOxOYL/VJxTq5KEMnCYXuAWyrwEUN/shmIt/CYjtRNxJXZnWkfhMhdC9
v7Y5v5iHFWCyIm+e5HUZKoUlJrA1qT5SUc2hkqjrIFSnCw4HCMC6LkLc3RVIJ3QeC/dhS9ZlG308
BD+W0zJYhSvMqNw0ucfNNaYoPaG3JtZN1ay5ApxgLhj1bKld1lKEyDBUpQt1tjh6GJIvNmwVGb+w
I2ZmH/TlBQNTt6NbgMr0ScdI/OtvNPPIyehAzWQHHbND/tKNNlQs+HUUNFppM2LFa66c1wpuk9w2
A1Yp8SPSoqBFOFffKiZ5acBnYDO0hEwm09QOWgaOzoHC/QQBqyoHvuNfxwmJzrj8gFccvqLaMs4y
r3ujZuH/MhmDP3j4uuCx0rke61Nm/bK7p3zRCZRURwtmVVQGxB9YRbPqHXzihcoUd8g5P95EGS1T
FfZ1dKmoY8Ewl42T7IIOGoqE1o6SLiK13Hp3HTlmXqediSi4yveMf/p1pQlVN4+IGDEk2eABZMfT
nRIrglPCqA5yjvJRwgxD67ZS58d6HYl/O/LQJl2ov8WC6Vcpr5jusItUBv9cLvyyQestv0XtwlB0
aYlyJLoXLln8fHYxiM+Wrb8btxcnepRcpLh/PjR1sx9Ix7ludAd4UbXeX+Ewro8ZMB8KdEYRIGQl
1Vzd66tdUE92thIBZBsYKKSatke5vtlbyktDETEQfsiTONvUiuafUjVNK5AwSnq2SLDBfftVCAiw
hsfFfyzk3iMQqpB6D1RJ0goX/7ihghhKsWvkq/EmG04lA5rIuEFRHcq7bxrDacs1RKrYgizq3EUn
oICQCH52dNEiYV2bXWgquHpmNsy3M2TOn+Ki4uiQA4lv2bQxhYAtzVN6muoE6OdZtQxEWjAtS1Xj
uLitXS0uPEHh2md7eaBKbkYrBYY2WhAWOMEgtGR/VxviwjKadON7gbPpKwQt7jN56i5LJLYEFdVm
nyzMxjh6A6LD9GDmXYv+Gea1x3NaimpGwIU0SvopyPeSEUoSvapxgyVjT+MmYY9nWT2cRqruYutm
PVB3l3rTk5PoPE4mfIYqGQ29c/V8tgbinnGCQ00o07cQMAHXAm+/Oa35qutpgBZ7Zg//qs0kDZ9k
et0rfaBG6X6SzGErlH/Rq368H+g5Z2fOa7fiDJEO+JfHpQvRR3dy+R7PXAq6G1Nkaj7NBYDnKk3Z
uLAa+ZRXjEpzYixJNF6bPPoEYp5TvsF5yfoH8IF5jBaDSBBbyBcgKJuFdSRrZ4KWTDIqcPJ5QT3z
XGortGGNZ7Kp9UjGVoM0sJkVosQER9ifafJDjh677Hy3AW31HloJOb3GNEd8GKDXvAfteUuSWhTw
ibmZRsf4NX14Y/dMAu455+gnQEIwNwQOttsM+bg72pl5Wg5USpUK4d/IcOErnWBc4oCVbFdALsoV
enA6l3xReV3DsZLf5Aa5b0vM8cmjV/nmlLHyLmyCMQUwACCw/FhFfv+hL3RI4etpi2Kenh5BjVZQ
H7yVJLhZoBbNsax6soCYH01z8MO3umXVXxYW9m2heeiXBr2J/0XkbUTx2fzQI+JkkeXZd+JPXdGR
9mBDgZszbFQqqiMPqEaxqiJV5XlCNnuOFStZNzBlCD/ubXDxxH5h3QxTAgmKV5SACfkzwu2UmLX6
kSBmipxfpnrVuDZUK5qEeZwThBdHgCuC7zQzQJABTsFMtJoEABAhsqA/GdPjIHKsrTEZ/cdRYG6M
9328+lJLmX6LZegFmTE0FN0ZCVVk69c4Qdn+RlXpTYzWMvJI9LQ7wx6ldtfkt12/PAoM0PsjqdcR
IeI8VZa8aiIKs4FCLUVAE7OJN955jBYT1VY9IJ2QFbefyIfM5UxondCgoi5uV5f1JX376ebX5ifx
ZZe2mWhDYeEhbsMBqo8Dhh0MtFbowC71LBTRnpciJGFq+0UBhtdaw7XBVcaVYDhxDI0rcvV4Go4X
TfG+4ZYRkq+IB+zcNhO3CXiFGIjXEbZy8E8Q+hyBv4DRglE1ncKqUZ1980aR5TjFi3KQ8s+hZazo
DZ5z70HDfi9lVxa8xZdEg2K/nSj9XjWJHIyNPGpYNc1IFW5YwBdGvtq+scRKdpdmHpj7V6ZT/dl1
jPn07v0pzD43C/RgHOsJiUq00Arlb9T0rsZhfsmPn6VTE7RxKq2rk+M01KcBwUV+pnLF0bDRUeHf
h7SWeNZv4LglxCkayxkR++tbSGCsl1zb9fCLOfLNHB5bt2GDZPZKInWfFRzUCP1h1AslchL6Qs+m
br9YnLkquaLNhJurViwxA7Oli+yOt6pL+1t8XgWZiwq1lL6HgrkTqZOrNfPwPWzVS4Fyg547qyhh
EFCyb5XmVKptK/emczGG1qLaUHF+3d6gw5lj5SCj5sRyRZKLD8Ch+MfnrTsQPndXjVZiQJLZaYZt
i0oLnCgVo7C4XnFN/G55rNZsw8LzmnUU2oVceHp3HW3mhV71O3o95nbU16uA0k+GAAdoZ/dzTmhq
Mr81vtggmvjvW2SUMaITA6DcGdRLGq2nhiW4giZNd5bt82BKNIzKPzUFxWUmvfbEXjjxj7obz/+Y
uKj2TfN1Q+/uePGsH0xmKXAM6zwm/rBJ7/wuVrer/H1cTAnX8EQc3AOQT6O17cXcYf3Hc7wMpCTE
kyoN0wiqZgzYVNEALNOIbYvccKC5NBfuL7vBDedcL2InFkzhmvXloJ/HtOAosj0Jmp67+l6LBM78
jgN4cCntAo6NUImXmT5jvGa5zJzeBMxfo3N25I7Rwauun/AWo7sKKjR/QyyAtWJNIecAHQuPYDpd
dad6OGx6chmnmSbjjdFRFxq3q/NP3/X+tOnfhcOgLBpMJdH6y2/YvbbnP2kgQg7ax1WkHYDaDIYQ
4oeDThU9docQJJIfAFNcFTZm0pAqNrSOFuHbbos6+fonZ9vg9GgcL5JEVKNxIZ+NjhygjJay0FU/
Oqe2EACX080zSOOisJv5bxS+MK7yKUwHAM/k5zwR3s7KZbr3nB6JKlpW4E54OBtCNjWJljnpT6CP
wsaDyJ3/8bKfz6yUBfrTYbHHB7D4HeLTt0crh/74mHRzHbO1lpo6zaxJFny9hIHxt0xewmkiKoRp
msZQg8eYRcUp5OctyS/fv1ohcsF04DTl/Zsz9PUM7y9eXo3vP7Ityy2F0I9TSIxzLmVeix+b0iKx
83qU9Szc1gsueGGVMayyjWbCOlwzHgTrUjKcAVyN7k+D/aeJbt9WiSnP32kKFVj7VgBiOw62LZwl
OfBmvR08Lm73nszuTZlzwYk4pcSkDUTmG6TRw+fKHHEfh06WAYQ0DkX2OSDORz/RXKJ3Fx+oIw9s
nfpmJ2N+HWKoBWwiviog6iWtLZ3UHN3y5UnoHfImq0j9aOkPJ7OGM8bLZvpYHz+CvnOuaKbP7gVi
JENcrHAP90WWuBrnjkKfNEjPRO/hIAVslxhc9Re+4aL3vmGzMCXHwvaOTtv6JXbaFeYvfUTKEEWU
63DtXddTt49EcfAW0FUzHuvQSMbPG1FCp3KvBcFMzOb1W5HXu37OornN8pV8EIMV5dmAkyC7a34D
V7niz1b4ODwVAzY39Uiv+Fc5Gz3fZYoV49WEzUBy6aprxdKaf2cl0IBFt9vu2S+0kXIZWvoWeDxN
2NABUCkNRMNqVV6fMmfIMt9COOSK07FZIHQJ50tTY6tXQGUxownzP0okLvHSmXGRCS4B1e+OuQKT
eoJtRJYqzy7omYQcgwUqdfYAU27SqMeTJPvr+XJe4AH4bPGmLdvVNBrPEMBtw7qWANwMm0GJfq7b
+cQdvVnpTsg6Xm+DeArL3Li2ZJE/2KfLCajZPdVw15MoeZUtSSHEeFT2S6Nb03ce1QXUsDAor6St
Q4hSRkT62H8Jh4yE1yxDPpg5iXWhT1Lv5DMxAZOsJNOlgKTLV3XDYP488Kjt5BATrGzLFOUMG5zq
gRagf1UetipBoqmneXujt7T18X3b93LZ1S2Q8DcnzBKFzKa9efMXZKUF47Rft1/qEafbaxbFjkuR
yQNg044QoG0ioczeIoFjVa5KVY0tB7XGjvv86YES9Ewsjfu7Fa+1qzGi9uwiwoA91TzAlqFwYHoN
XFAnLKf0MWbDpenrXTS4DqHPuJQok8fXWPUte26yhvIFjR5yGoNZJ4Ka70lcJI1AHfedWJCMBROH
/cqcLv/tfn42IpgzHZvfyfzlopz2dxZ0aSUzNjkd+EgrGu1VxLtCao+0eQQFtzc4EIO4x9U73Jfc
AVIhxBaIscyef5HX0FlCpMh5Fg8DoXPVeHAEnwOE8/iuapAyxEUOEyyxQbJOGrR0MFg6arvByQLy
WF0Og+T4CyFZMwaiMmvPf1/RQqcypfquQ9jqhDWd3x3SGe9aq+33ZZI1xLIKukz9an/jqH4fOKyX
T+f/7kslQB2nYVXZiHlkRTmAYpqGtME8MO5iL3H4Xu7x5aIl/iixgok6uZuC9tQJTY8Y9eG0Cba2
M5ctQ2MtkwzQ3tCKlbXTs91koxNYtj4jVliKwVNxcvlKAwHQisRyvU3ikhq4bHBwDVXzRQfPSTgs
KFXIwfobeTiuOW9KJ92cqWJouT9xKTi2lu2IzsBtxQ2AZLZVwMPw1Sv2Ntr+ZpJeE/ExBI3AHtw1
KBv5ji5GhaT7V1b/ZuM6wgdLufMCne4aqfr/89KqU8lVy5JPtUHd6xbM0UXCXUVPvXV6QD/LNUL6
ZChFOqVgogGgtHwXwbKuMC59kf54L7zo0uKlBIRfE/+xdQMaNz00ZmvsruAOc+keIGvZEqK7/gOb
1jADiqI8mTQrTIgBwvFZf+TaFx/BhOLQGxl+U4zh6Ks/khKB2cuMDFWb/2OgH0LiS6OOLSrwK2zG
VEFp0ESz4hLbZTAt0HLnFt6+nHCkjo1cP7uDX7BKsYF+j9HBmh0ZRRPv8pJXecnF+ozQt3JSZ91m
w6jl0tHI6yPlAedWPjpTjsU5l/KclNZxx34050La14r8McgpWC/kRWwyrW/LriWvD0VROOs9Fvf4
PyGddoRXCowfbLvFADUSIOJgtlVmlN46pZAPEVbzKK/XVvYt7NGOozw7GeAIEvmqdLVjU+nElQPS
e5Kc3jg+37nlNrEa6BWYULrZPqxkxyZ4wiWVDuu0j0hDlt+llcY9Y16RencPoyrlQ2OT78wWzI5J
v+8hUoA0FwBsyqsbP2ovmUZtFrgNdYDh/inf3MDDETvA6D7vLE6qpySynAlpeNDkF8F3HHRMPbyk
wqSYkMBwj8/bFPm/9UqSuwJ6dNmBz7EWI8gvdmBlcAtQKK3oIDc8W/061Lw1Aa8+SGePtqyunCBn
NWV6DPBQf78SalMqpMgZ9MnBnGqO+LPsG2WUjQrAtaF4iI+2Lt4cvAw6dF5LK442Zwz+f8T6S/22
ela81w8OVhpDF4byxvsgr4SASJ2yau1lRugmyPKDO+h4o3bUICQcywzu1IVcZDjM6SZguYS4WbgG
KmX9cC8bV4ayj9QltMClNL9wrYl3wwn+mAPSFIbrze+HyFq9y9mLxIDlVEm8uIOGAjDA6JAYsrG6
p4CSre3c6w9lerNPQp88GyWQG4zdYDG5/SOFKblNl6ada+eF++eG/oldkdEi1Ww85cKCWlppt20y
wC1OlKuMFUIjOSRG7YmPF2nxWoBg4ECsrxio4fyE6pr3XjG6cxkl2gsAnHohDRu9UTQsfEvAeByd
qtHTTrvdPCgyqdK9ejql+zvSjXG7pyNCu/L6eMdZnSntucYCuiiZSDGsRgcxgm91eYuPYdY9i88X
etnlhqkUsVihOyDdouFIlkLcoommr2DtJBd+/+lfF+aXGYGlZw6vo9LZaQcJ/tH486Xvow2PPQb/
5tQHrcNSwMJoB9QUnS6cOUyywP8co4ETtyk+jQjwKu9wp1R26WxjygLwbQLP/F1zS0K8DzCdRh+u
4TL5N5Abzf9wcWf6ppfD/iKJN29lVIFRjjh4nouqoHGIRruhusk7r98LaH9EID5CrbztwxuiihSv
KtKYCRGkoiKC1OiBsE/sVeRZxPmXYvb5RNcZWdlknzTi2tWG/T+AL1JclRopmEbahCE3dGjOYyP1
eDMe2TfpQejwvY/tYXuarLXMsgvTallaaeze8RTJXXHAmzcByR5I8DOAU4jTEcdEtNOVvl0z3eie
DY21ukJjpe8cf1Lyx/hEsfMsO0D/wzY/EO9f3qM8DjkO+io9GmcuNpW59XTf7M7tPqLcYj2q0kPb
DA+G3EgXAHgXDtXCPitkwSM8unzpGRs3fWBlwZEIh3bUcCpyPD8yNQhHSln9aUmZepUyPoYD5wxF
HC+3g/BWE0SZENdkJt2cuyumukOlwFI6tls5JSyPuOPRtb4ZqcDwAvx4THZVlBgq5EGW/z3+b4+V
TyuEAbMV114MoPaQG6Ml8JgGZ85GRk9ZMyHFyjK+//65MkmZ83SkE4pQM1wOBvh7NzJWsvmhC2fn
2MauwiMjQOHLaprheQpp76rwS/+9PA/qZH3m/ORA3/MO2+AASZT4YcWZ9iszeoo8HIHzZP2EliRq
Aq82vTA9J3wjzv+UZIv9uc4XhUkjaf90wctcqLc/Tn3D9cJ7pNtHgnVQ7GzqKl1dSmqSKUiYeBQh
5JbUzTFca9ODQ2RQdKhh/QIAN7IaYww3aOf/WyILL4Ut6LfJDgI6h8BcVKrsdh/AQoAEmQ1tC3Kb
2qPhOgwtepLjViwf1p7gu7ZrKVd2zDvFJiVh1JRt8JEYT3rx5bMmxAc8gM26gVMBv/2RS1xpZE8e
5E26EM9OrOzs0P1qRMDZ+CLzlLlxeXicx4qtQzzvAw+Zz7oa0WEIZStlCL/KmF6l0yUXRxFH7PEf
ie+FMWztceXpmdUHs6KSLpdfIL1WRajjU8TRWExbljkjMxuoIRwnfKDewq/UuSutHa8Tri3v4r8g
ZgZ6eoHPey4/WVkP8CwNzvvDwmZxOEW6mZ9daN8LfKN63g3n04O5AgnHSkibqo5YhNHKQce1nNvc
ZvAAz/tAfOqSquX7ctRa0NceHWnD0PWs4vwCIagq9KxUlBOCl8jWIJBUD8ElOEU2Ec9Ftv1oZKWP
hIoa7gk70SrDPS6BbVLvE09f82TfJynRftKTaQZvUCpdGXdG/kpgYq26mZVsTdoJKyAZPp/IpnI5
grGVGKaKhZODyO8XrtVzFNZAkno9u6sK2c1yBngdG2Tm3ikCUtd80Op0NJrFCthscdpDWB1WBWwg
HG40imEb1ong5pKyV3ZZQRzgZ5REIuwhXpRITOzhprFsXfD/ZtTzR1MH1ik0SYp1pPKXB2RZ+/8u
bgBXL1Zxow8Wdlsv5KsphljfHF+TcUoBeEhSja0DvCPVpnilidTkysao9CNioDGSsmrKC3hVkJlh
2wRUEj3FJwOpWOLP8/KnfSyG55T//FHpGNDIYdR1CCrZWwlqj27lo7uqHWVdL4QYsimxyFbzn3JG
0VE5t6Ce5KrelZ+IUIelF+4BIYvPAMn0w0tCWC9BM+FkD+gVBZmqW1bfFOjp443GdYdFtM9AkE2J
gnKkaE+nGbpqDY8d5O55rqJUmAJxEZrkCN3iq/sHiSNZxvBZGefGS2Z5lU86Rl1Erw2R7/xuUdUo
le5OrwBuG2VOiOj3Qfk47HkLnn7lnFVWdcD5+HSx84x3+OuHmOePnexsCAE10Vkos2KuTzLrQc0S
t+zwYMnfJKubLuIe6eVyDs/s/5EacO10XNEQuUTXBLmUiOyH7/7ibBN8mxkeowZwGn5vkk/LYAN5
gfUblurA/FlbVIro6UAp2YZYmAwnKZC4Y5svTxpBZjUMW7gH+aidhhn7O2BKdxjAqD5wj9pLOteQ
QDB+v0kD5fmkFQSCaeVO9helQ4coHlxjztrAwVxUqH+g7ph4ywWjH1lidJB+IhifzLMOmVrMZlvj
Ixm7sJaWq2SBJwpAAkkDHMMgmGEcDNSpNh+0476QD0AsraQPyEKM20ace6Lx9jKUQIqrjQ9xKeAo
ulyGQ2vv1SKR7X1+Ye4tcLtc55P6hElUaYAyv8jV/YMmJfCKydcArmzg/6D+v19EhFIwTmUiSV4o
EjK7iW8MyCfyTozW+By1fII0CFkbriesAjGNcgSifmnoM/vp6tmRdGwBsZdfq9oUebSQign+CrOT
GukPqkXM3uqfKmJ0xDYMbAcWPCtXLFWLl1qgzFdF58qul84BqL/4ZRqmD39ZyxT8+EpafY6dWo99
JXcbHtivL14j27d57yzizgijAJkGtEFUkBA5cta5dRe054Uxd1NjpaAegIjIgq6ppDCkM5/4SnQ5
AMEqXPhJ4iqMLWmpI4QnVxuNA3BN4rN3rAMF/Ko9ipV8ffV08De8vBd2SZUJzpcxYn61Hufyi6i4
MAd+mS/5NvJCshqXsu7ToGAmVKBuh4u4aMyjgYoF/yP1uOikrMfgrTuA5cDTgwvKTdtFt2ucPzMT
Ce6gGPg5aBBIh3Yii/c0b/+GgscrZu/ru0p5jZCOCLy0VtXdI1hN1JZNF2qvI5X0UVsos0zE+bla
/oea2nUErD2awylZ3l4pzkqA6z14G0Y1/2w1h10bk3xK8h2YrogurDzlbXHT+F5viKmlOyOzr34G
9KB9TqaidOyeaeSIr60vcmRlOLWqRMaFn7M9k0CPh7WF55E28A8BzCt+QKRWAIwW0+iYob/SlFS+
rvs1Zqi0hRXsOqcLCE9enu/tnknm0sAejuFJWqn7kNU804S/uPH9zgjXXfLfB8SUtEkwraxVt+oT
lK4BJusZi5a9+5i7jC4ipNYQfqp2aRLW48RtTR77U4jKd35+aMi8gylEzMOrxsNNDN4WM6Rg6PwP
kszmLsG7oNKoU3+1eQMELVRq5kJTDgTJEzyOi5As3E4yH6VWUD+YHdObCVYcS+fuM3GPCHnKllUw
CLMMvcxbixpA2z/ZRtx1oI73Wk+Yl35L/xfYiw5FbGkZvBdm146HYgTkqzbkv7Qywkt8evC5mMqX
cpV/NestYwJ5vyBqm/6UsbGbqoWWY6qKYrINU6kmRL6zvXv3DLFbaeRtxD3g10CQG6b6aYOTwpLa
fT3NH+yg+SQQUl67deBjdxFXRKX3fs+O0uGeIRWbkwtYaAcg1kPtFso45WLU23imIA1dxAd6oveo
hmsF5zCGKMMxETV0syiDeExUXAqLRjoUfjqVgczh1TwOKEsSXp04Ju2Mq8o1mBRhiFMkQIkdVTKc
OVoLcVuQrQhpyLWtrue2cmCuGCr7w9PWgDfULDwnJGycx4MwgADn7pRRYzfrouLu/hZDqYInBd9V
5EopnvrDdDasSP8ZpiIUHoFlYA+1Zs7DcZE3by/jGJH9+FMer9bSeSxPBQMlu3qdhiyd8en/8Ocj
L/OCyHDBPBqgqQK9anekt4Ro4cndo7VL41c9MnbdZ0tnPJ1NeH7DCmOBKA+lW5/prCKvHtDAI9E8
zYF6ovwnzllIoYu4wmMfLE7Muu+LSSx0Qc4NKzfnDiYSpbFy/MiGfIaNRgGA2Fck9jU1srLxdmIU
4JZHdsou8AqWY8aBmiqGfrNNkhLaZt1M9JwbDByGg3ltcmcP/IoVKuoGde+XpkgjslZ3q4SLkDsk
yjOvWl+ZYrrJWrI27X3zUQZi9qKT/blrxVJ9mt+g9K1juG4I/J0yyD052cSBZe25uyx3as9cpJXC
jbT8u92/m27f4sWyNZhx7bAy7LrloDQ2ANVWGSePLTxibmFwYILaTJaecrYHS36lgCJUu04TiF4P
gYp3qo6UZw5iVVn1FmnGheJIKAWc1keOSp/2r33S18BG8MtR4VdiKycn9G9gvOKDajVa3c2+4TPd
LwUjKGQ0S8ETihd6SP8F0nb+7fKDeuwf5z0QsaBRold8b7T22OEeD/4/waQVnj/5cs82fYbW9OLX
1dSVVZBnJzUutcf8TAXz2W/i4sxTkM3A2Cg1nQUWyLmLGlsWEiMyvo0mJs/nTLC4ZdqBTKJTOgmL
9imckZ+scd4d6JKNpkWsuqXuMw6bIbfA6AoMGSUm+U08bMl6+a826bNWcvjPmvUL1Q2qX/MKBFE+
S5rO4MjJiyMBqjjyeYUNXBQfQo1zjTU9WmTvfBi1s/jREK8KYU4VseFSu/bZeEfTi1iKR7FmKws6
f/JZ+wKvNL8Z++yTvEX4TkTvYL6l/vutJQi6UebUCLyR8XzTFQI1Brnm6yVpQ5mrySsVeHv6tosL
v/BfxWAYjZzr0/JcdkI/bdrkIiQSO4ovgRIaPu4tR6RMV/HuQrJpOgxvbmpHmQ3SREic65RNc6mN
KPMRsPLS2wHoVoJh/s/tLTACUrnRQXFppVciSl2fRqKZi+qNFf68VrKHMcVjd7dMqxrC31MJ4oMV
xIMswZAKuC6BoKxOcytWrc0/GUw30fqS7SNhvHAtfR7K7zmhjjezDghkKlT2EXFn5xH9qZpvIVQR
IQJeKSXxlhDtv2rI5M4jaRiWJ25OjH+rZfmsiS3FKw3GZiVPkFSk+cyyy9fPhbSv2/UmK2X3KWWT
eONxTVR/rdoGfb7Ox4sgZzrs7WKWiKNSOl2N2oR0gSEI88geFA1GiPJah6OkgDbukuNXabexHv6L
+up+JWCwkCa1wMJGbgP7VpZXII6aDLynj1alD6HBqsDPP/qty1iJ55Y3kfbfpwy8XFsoLPes8nzo
Z3NUq95/r167PNnvuF4rZQx6w93DjKhLU0dRySmtqmyjI9hldlp6KSj7QkUVABhtQzftJDr6/tV5
b1rYtcSc9VWOHPoaNCOyI8gb2FWDQJcUYdsC+nNGT1yX6TPW7lzr81RLxfu44Drfjt+0YjgQ/PQF
/d1NVmykeZPzTCi1WrOOjeQVZWr604abKMOOy/nZkXKswrHgDfi3jeRz/J3QP6e9KRLQQiIboRgD
xeNqjSrgIteakX4ckj4SwfoJ4KWyBiSLmUTWtnI6IES2pV+oGSc2w7BmRLbySNsSCKGDueTqAfLC
M/VTKNATWHVDeK9CtX+h8vkamOd2PX5E1oOi22qFP7zAtLDFPI2FDXMXcAUvThRORGMs/l1Bd3Q1
58ZMmWqDwl9ctimiNuzPVKMKugEmh1hDXgdvwQLGBXIMHk+B2ArksHeOt6z7qw2Yhf66hOKfYIb7
tKMazEpmN2ON01PjYTTnBaNpUrWJJmSX6z+yYz3mEcLDMjeDSqO4BeBoXl/qBSIyAwQPTl37gLhe
2UkF2SAvAwqKstQxQEgMCJ8xL5zp3OoBAu1xgTZMkVc99F7PvWC9j7OvvTajv7cljcIWpf44vioC
dFA2sAEnkChlG8h+ZUbD+hK3+LHqQX5/9KQhNkkWYQjJMAKxC+ycuo2jQPTklKRtxXeS8zzqw+PZ
AsxkDUK8LzpA9ANUas2SwOHUndLcOpHZzrdqMyRyrVhn/Em3DdXtPvLgLtAyGFKjTirqIeoaFnKI
5jdYYIy/u28gHkk8ZXafxftVYgR+3ZLXn9JgLg0ISyUdpXC2QvYAnxsPFb26/Au8livltY6kzIqI
mwDQeMmvUvqs18U3T3P9kN/yvJKRw4e/7Xmh9nNJSy1NUVjA+1tyWSrLnsNItAfwiuz/vQqPzcob
B7aJY0K/XArdOsrnUlOodqbR3+cKVjIIu4PcCjsQt0MtZIWUmRraVeanSznjha9pbFVJCscaLpn4
X0/ii5+Zt0sybaRcCOVVuqfvZoB1l4aQF4xV1H7cYzzcza+F+itgsaknN2aWdIlHlQBgT1L9s6mj
pDJNW6rvjtV/qFT+9zX3+kutPvXDZaJdll5UiD1YiWrXmPUNpfOU7QwAjA7aoY8YJUxCBQ+GtyVP
WufgDvcb5hk8w2oRgdZZb7oxtYNi6r9YebrTXLPC1XBM0gvJCVEXUCVVbgtI83CK3CnperAzQaE+
C9eTWwWMzaVh9beLOq7dIvCBR6Dh5Y6OjDgTfTW9S6Vxpk7SYwDjVPNb+wlJ/Bz4cczhR1VrWPf3
Z4oBJDABQBe6CQwjGVb7sAgdXjiq6xGSV3r9QWmMOFNGrKcCYuYWRWkBTzL+zlKDIiK1Yem8LEHX
/pMzBeR7tnAZQxrqpFKephZ1FDwrg68wRE/X9DBRCgd2JxJXaRepD80WkNFjj1UgxH46vNxUfWaG
WdbNhsaLznXUevNOM/BZr5b2+9bxDlEp/7MWkBW2ZTy8pvpI2RBxiD/kKlvN+oVT8F6OK5pFvIbL
DI/K649W0ZTVRGIf9oGOQe1Zok1d329ifE+iyd9+GuXAmlqvh5KtMEZwjWJtBNzsfCsz0dF7IQeU
P2uMAH0Gf79EkX9yZPwWaAkGaZLkc+fhEKSwsf+9Bk63xqU4mH4EHQ4XZCNeB+4uIxJqWefKIy7e
juQ/WVvofB3GylHEiP4YTZCieaco3JVSj7sWSFQQiD8Qa5IKkDQSDLwKhJK9ho3CFpZiyIakZdIS
wNdCoD8HvppFNxPmX7/NSy42YwluwreGzNWsp9QwPgYjTNJgPT3vPyoBL+YLQ3VOeWOxNTS5Zhq7
bkn4tvYLzzVcFLwY/7WnTWjlFgGBBVocYKTHErzwKQYhYmRC5cpBbxP0jm8hnuOPFEVpsUSXfm8v
SM0mWd6BVQon3fyrU21Eb3Dj29UiZ/zaKsMlSL/pQ34havFezlUZIuw/Jn0tRvmN0SV8ezo0c/wT
io96mwofyV3w+SLbePk0SbeL+DekvDk3t6j/ODNsApfFEX42gplMWTx9WWCFSmlydL74B20xg0y/
PnGC+2euyd/nIhuw8P7e3QKfQoGaA+kleGjz1LpRevW6w/Z6VMGSlDuWEjLq4RhcFQKFGt94L0L/
5cCXb+53G+MlxWkPbY7oSkSsxNnYGQEKbZHZ71W9RyC8gEQUUOL5VxHIG8GYCGOA6rSLJBOa6Cae
r872zIGr7Uyl0Zf0CCImuPOdx5v9d2hnxSoa7RKKtCOzV3703OGaekBncctYk6Xxt+MgXEskV7j3
Ydy+b+GECKZiruHwKPxS4V66x/0PZxhluJ6W6siSMAvt0rZUBMZbsTnIRZkrzPlKY/AJxObkMCw8
ujX0eKJVlyADVG7ym1HPSktJfkr1ir17UxwF7il9HXNOV5fhdJqbwTvPPu7Mm054+SGtVM+gilnC
wwWT/oUVT0UIr8u84F4AunuqVp8EOWwSvc/iC7TaKJXlhy1Uv/Wox0kJzJYGvDBN6D7O/m3U1Zuv
aOcXqiGOQbAW9jKeOhbH+/NymsHtcLscPjchrToVgUBqSZwFIa3FXxAzbcWBvxvCgqXyQnrl5//z
hsdv5yBrUM64fadB/Rb0L9F9fNkw/gQEOu/r/v9cHs4QzKp4cmBqf/AuLYQCEb5A47Zd2Yw8iGrb
ow9rRc49pZGVZhxcKDSepHfqxjzHXMidpskXKJZMEzqRbKNKHJEu10yBAdyNiGVfMknpXD0iNowT
e7KjB9BrAflc/IHieNEeJw/mPv80Eee1J2+nuFVnFabQIUvHIoVNv+oGhzhv1EmtubYPYiTn5g5b
OrlQRKSlpaklpJNNQ+/iu+0M9PprBuLpf9K6XxdDd779f5CZqmz88QTdzEJ7vMX5mDHT+r7e21wT
e9EebkhQ9u23Gty62mgphdnREAvi4MxpkjDX/6sgHeUKrkqlM3hAQOmWHSZMSNWD994d5tSNaSft
NHiL/PK8QXhvD/Elc9uhOClVJtWMp9Yz4yUuPjwya/14TxHisY8hZAasH2elqdGocVAmJDqTZtLK
hmFAfG6OulicaVb/+8pkpnjTKr4yNnM724fFNmAotINwws9gm/tH+0kT4tdqEqPV2ax3xFnBPIgs
n6xvnayp4xSoQVBIX9MSs6xQWuQ326kkCn2IpLBCovBiRe+mcxDffqmDaz8Pmxr0JGoYTbyjaZjL
GWfx09QD+JRQpW1qKEfF1NJWp8JpSLJVt1phWEcbM4Lqz84sBEdBNmtyGZ4mfIayfdPXHLu8rOZw
vuZ/jPnjQL33sDQsYi2lO6/+J9Tl/aUmJGqYPgWkJuwiz9P3MCKWENO2ZkTuG9XQxEiynNcHN3lb
WWR4HtVJMGprL92aLLseX4beNdnGulVvFn4zfS4ByP+CWNoGkR4BRY0jg+xI2ORTj1AjbRBSsXaF
WDWIHgcv1tTzNTWzmrFRpA3D0NP0j/sJo+z3PjP5Q6IIho52nhqTCAJrk1g4JG3Fc46jpXz0tlpz
hysR08jjbpcW5kQu+/ohgBWygg6qpF25u7ox8MFVtXyAm0bRZk45ARDtDPHXivmTyhVHx/DqFdAB
jwLw+rbnOFt7xvLZTvFMkYo0BCABX5ncBwgVeB2FNhni8EZwFGg2BxkZDnpMXHv+ioG0+yzBf6zo
6mjJsZNkf68r+oydntO+JoPQRCOKK53bMAmrRdY/ccekEs8TtT4bWyFr4iboDkESfgQE83JlHj9d
29Vj/FF9bLbyl0HGl+qvMdID5QlMJpALOD/fNFh+UsB1e/zloPisAxqWa+toBC+Ooc37ZrM/M37C
wUoVfh+yD2HvhDJPAKHbrcqVpYboNyaWklnTDT8FtYCbQBgaf9mlwrJa1CeV1ZQ4hKq4j07PpFOT
tcsZAd6PF1Y018LwvdQX2Wp+DWOvxzqrRrP18c55y5QdDg581pU3OsQInTezUUStE/yxXqXkBZB8
n4SPw9tCIri37O0ohvlHuYgvwFEJUH+p8i1+QwOyXgZ/+e9uER9KDVpLsUu+Tnxc7rEwO7nJkMRs
gso6mXnCTngx7I0iLYs5O/zTwqQ97+fRWi36bge575S8pdJ/Pgkt8hqjlae+tViGXsVQV3ORyEyI
81IaUQaI1b4+eiaFkl2cktTtbNwHsiHDzDjGFENFuO3pWSm8NnhxvsvjsOngG3DiTz+0UcN7yQ1W
goL6mplVerYApeitLJ6t+OVy1A/zJgrTvRZcXcYhhgrRl2j0u8808kUVrnj5yuP63FDpdIUlatku
Fwr0Mzveq0seWXij5TsFxbV1x4enOYB8z9AskU/EoyEusuUxUJfGlJanBHf+KFX3XGrdfCX4jr7M
Qv6TvLsrMyTAN2VWj+Mt3ETAD72QjY/55LRbQ8Lgmn/yTPDOtOk9z7wWQprQBd+nt/Gp59H/yo+y
eC0V/9sYSOWI1M0Ki/ExsrLdrIP/0gW6Gy4K2O/l8s+TfkGVKUsfSnm3LHz1wRVKLGI65CNj8NxV
PVAi++BFNbbxTMw09i/WrpYCleB2o7YFitBj++gVUEOv69yzKAgcewQ2N5E4bnunG352RcJPLiL/
blQ45uFCtuhmCp/7QeKjy3fBfAMNnnLLACnTaUHRzgLRTLWoUdyBGvpg8V7YHGB2mnM5KH6osvIU
wzJyDJznVZJTwQGuWvwnwObyiWrOHdRLpwfk9pERqP3MpoTGTK2zXarf3pWT9L/tx9uVKCnM3uP1
gT4sYfkGoOWl0Z0LdScYaujdZ91J3LnX4yLpslMenAXw2faUMf9DpB3gCtPHggfxMhlemPxxL1KK
ZimwTdpbjckV3D+9TJN9zYfy3uycg1xNxtnO9My518WBzI0J8RtbXSJodT4qlDEuihLVqoLO9Owd
bBcdISiqyDMYL/8FWE5fszONOxzgIDdSV+hOxJIR8T6JLHcLLBrDxRiWFnDEwxlgXGKgyA/B1cjb
0z8fl++qqPhxCHyzQYiPKQICoz3cRdHrFcu5/GNKwmCI7WrSDCilREXXP+YEAPUJk3ZHoO5jjsM/
ru4BwYwb8wii9Xc+v2FQV/MCekCWt0zx/K33e4y5qsZkLOrnsw0MzbK8i2PH/jg2MvCU1OTDhwai
8rkSEATeNX5CPxB4jfr4+hQBrxcUg+j3o0CgjbDqo0KQcISRQmzXyzRUeFMih0sCY/PPBVVgV81X
KT32z8oaIrfT5p6gq1tHkQ5wLV+r54+KJt8j+hzYiH4Ui4JRzOfeLSKjIscqAaf63guvBznucWlf
9wfIF0hfMXu+bXNLy6lK920zCpYY18cJb/bPhLdbsMPmI5pNJ7T+tRWZvTGbMjcy6YbeIuHj/SQY
pEbkIJBIu89xC5DH3FT5vuu1EQgceFhS0wY4mgMTi/rqSYntv+m2LWoi3QHe4BvV/gJTKxp1ZyB6
gEYzvX4INmdUxUHlNBREu8Q+pWBec4fqf4xuAEb1J7a9UJ5IzIGTjMdfp9f6LredAAlM/jvSuyPC
O8MooFbYy6Q9BcF4QLsq56XtJGDWM3MT341X+3M1WI3qFwMt1o3H2r1Y5ta5UdxfmPNfDITSLuCy
IrVYrXumyHKUXUnX9gFdW8kbSvKv9K6ouYSHGCSHW1UT8f9T5kGJdORfCU7FLckJ+SoWLZmZuu2J
vVEO04VQ/i1sc4kiBMsi5fsnaB/xJQfekA4Go3oDqISDKT9JV7L7rVRHK6ykKS90O+3MRw/T4rRI
MhBeRakg+4JwZ8C/tnKKS5BDpHk856n5P3XcCcx3dxOImcepRzi203SoDruCfuvMimVMPER4tNj8
l1WVLDH3+rgGoXHk+lWbeihwfikpAQCxlft8GooHSHw9xVKHVEjV8HFJaEuAaJRT+n12YhGdwxgh
QU3HILsF7zj9dVgDQsMdiwI8DwKEv/3BSGt29+N5a+1BrwfoNaUN093pAv/Z222Q8whbniDxSQVG
Xkw9HSXDzrc0PzaIGjhsFzTwYvD1HOevsojX473bpJwV6qDinnnBqV/Ek/sNv6SWhM4sDnDkecjR
2U2jrBhQS0EsDymWbn6wN5XwAHSv/gwLFLUdvy67Xcrs07uvTPbWNpqOLuHbxcBb+dd5MU6qnV/R
usVdD6gKuaM7h+Z+bhSxoseifvbOdL/NZ0WSI0l3N04q1rhpZgaVQ9voYsoCZUKJ2NVIFJ1vhK0L
SsZoj9+9TIJ9OMEH8ZqjrtA4fBn1E9kWVzFRohHsux830IC7/R8rfwldDkvViOzl/OwHrkRVStNf
yfdgV1kmgk6YFUHjnjY1Bja4fnbAEWVE1iP5WzAKcETgXkt+ZhGu49s9o4grSbYIaVYDmNLU+rpY
2exCkG+R5xdcHo2GRL7rIEtMuTDxhAphyI6oWVw0pRrkt8CnlkVIjS94ZjfxEn2omgHV+c1Mg+zH
kJsFVdtcn91t4uqV8ftavGGyf5Mpj53dhL28eNHHARmd6uIwYFicp4hL/zjeT4dEg/NOnTzndQcv
Knv7WqKwcLEMRd8wVDJkx1kLG5Eu3h9d/DfFl3qZanq/toQNdTHd7zSL501kOqMp87xUd7oYN+2m
8Ic3wZ9dOm5Ftv7yHsurBgp6XSjoSuMWbCK7GVEFpxX4rOQ1zLAYd17FrinJo9eYl9sZOgmfmC5s
m3qq+lZ5T4M8YRzFiOX2iL/QSjJpstiLOTIczwKZDViKiZVCZn4ngRg0tMe0zoRv8xzaPrqaVMpQ
N8wfYR1MCr1pOUOtEHbNKSKK8hHKOV/GG/vRc7JAg0Nm0FljEzs1CJAwYmhn4LlPNM70E19GFiEK
PeEkK3VspkROhYaHas35qG4zYdJHEqQHdoBeC56GPEQxPeRmpkYOHW/QqIvF9ESlhADPZZllaEs3
0OH7SDGEIJap0/Anhz58fTFw1gCrBO9uEDDitM7/Dbre+npgznlWIeu83JPL286Opq0Ik/mkRmYV
mhma6ZtkGqLMwDB70m9hS0L+4DgPyT+ZeRSd39L797IY0FV4qH1xtwW5oc+Rn7tlZiZdLyCgQDmk
XKuIw+Mr2StdycDdzEQzT4CBsDDDnU7EJpepQcFPgkyb0IsjubrhSiJ37Bs2mSPXwHMHNgC7R+06
81r3CJlFM4EE8F6OMp4WdBb4MUNsWMF/ydqHqIZ7s6tjI/CS6uWle2xFSy0KB6cNi7wxFaP9zSJ1
n459AXL5lrXw/VtE6mk0GcIdyt5JqXWQzkc1oEWMl1yJWrzQC+VEWPuQEQG6tDxAOCiMlMOza2mo
O6MPcbRHV2/nkPX9QsO3PkcGl8NQnf0MqVz0J9qXZzA3AE9FQAdiyJRf73Oy+HIN7WIdHOPPY5lt
yVsgnLQGTbondUQKkUvZ5jbaXMEyFRyPMe9QT3jXr72q86xkrtc9+3fCJqri7FNvm7g5PmzK2QvL
AlwuUSx83qzpQQ+bjFQrzeQdyOrjjYvWcDwu9zm+J02HhjVzHd3857iLjpDveHg45vMJKo7Di220
KbF3/EE+NNVqC206rglnjlIrIdJLs+nYyJXpSe6U8u7r6EbdfpQCFPW2yCt0/6iJWrBCkWKw7iAq
0/w0EzaxjeksT3iuVxqBDCg0oyAaAHtK25WlqcTwPfObLFnZyelFfi6H7DCMz0q131wd80HYFnNy
0jJlG14pj0ncdHlM/RG1VBtiLul9dh5BCcoVQAQMu2F1SeNe/OBXy86afVE+E+l0PgdSo7hfQawA
vhrZcHUpulB3nVoxAdfhVfpha1e0oAChqk02C23f0yme+FSIO8rHsIZw4GoY7kRINLR2JVFUy6iF
VxpJajoPkLIdO0ATR9ZAYA1RXxPCROnqBR80k4UPRkGeUCF4GYt1oMbybS0hqX6xV20/AVTLLOeG
l+TAEeLdLJwnMyp6NCrnGdYiVotX8JExKBG8uc1cVOkWrRj3anVEjJcXNdda+6o6Ay2j3S0OGnjS
QKNayrePZ/71+meu+3eRmlJsduCCEPMPuvYMqISvAelmEQtGbNSmmWQmm6lhbAf61Ar6M06jNec+
1ypfMKEt48zcq64wUxF+86GhXJyuo7sOCku1RoZlK80FBge9mEjrx5UJkPwRItBxYoyfj3txtbJK
A2fhoMAfdHM8NmORWo/HGmz04uNioARbgtbBqtr1Xp3RVDSMDhfM8wZ3HlXz2t60iPrakl7PNIIN
3zuhCRxPvwTXD+Q8w9wi7peR8ZiXJqT+E12D7HxKHxznkuHBEBcFdvrvNHhC23NOmksvee8VqURp
AQ5DwBwVKr91CNu0jCG6WNAJHpaB+L0wvuffJZ8SjNZlVg/V2nLmdzN7+TzUS44u1vGiW9xXbcKh
wa+htvdh2GIpGiXsrH+bELYNcm3xnzdPJEfGAIywkHawJ5xPGap+n41TiYg6wYYSqsQCVjvBQk0A
gMRDTwO7g+sWfr3AacsyxJxs9yhm/n7N0DbFHNOg3C/74ts3aQ7oASirgH0EZfD7UYL9379VzTCG
GJhOqEs0z9d2MQCzxr1AYHgiG0e+e5btp/3DVrwluLQ6gWlZKy5W4TGzWadspEwyJTYF40IZ2PBJ
7OlzEahFyMy4BElqlpkZJMVktpCIPQJe6mzymI/5w8SAV6v0Fyv+M9B3lTeTEC7JawNFxSQBnJad
KcNxytuHKv2y55FW/Tb1205uDLPYLoxreXE7jaeaX/2vnKGx/vai6Xot/9os6kguVoYugvpV/tOL
1bMFr9gu0d9ZcAeZAcPPAk9GoS44Qcn9ZHT7gMLCpSkjDp/Aq5zGvO8KpTB2TIDbwvDdrIlSBYa5
0NSKGgBbYUsqdg/W1BUEpPb2lea3jOzLUWst90ER8FT4ve7YCoCv95IJTmhVhs5BuJWT0MLxLiIe
KKMg53g1vU1KToi8l9nu6l5QMvCpfN+f/NjMNIutKROpPmT/4IGwC77TkAihlVVhU5VwJl6DXluM
9bKMWxbDliwdLPAp3YEUCa3vPWxANG9WysUP6MMjGK31BBXOQpCusflNqzso95Lhfrk1azm6GzJ2
TYC9/eYvc1HUCigTlbnl9ePGWDMgcqqAf97a3upnQGZXx+CN+hc3ujfx56DCcwwjq3FJKgl7ewbA
Ur3zkgvvMLnkEZI6I+RRrdfnOWa9RNXIh7aQYx6lBqFw0pS2N4yPTsgmHlQSu4pjcDrngM5GLfnc
EAzLSSBeysyrItg/C+3WyTylGlIr6N72bLKhIaReqpmqnNCiVU1J6lrsUCTLrxy1Aj+QgHswFZLc
Isk+LpvztlVa/BD1hOgCOPHpP+1P7sEFjmoBJjIPrvNo6ajAWMnE10aXo1oZpYKNWSjvh/9UMfjz
2SG2ZsZEKXLqOcDpbLyqn1QGqqx8vucMmYrgxT20aV4KEDEYvYMNuhh4HsRfPX5ex7UtyuV2qYPx
wfyv5tFEKAkM3SRdTsmJIjRLHZt9euHUWOihk6MaZX68wdqa8yM7vArlbb3+7yi3PO5ErIVBGUdv
gqvclbXssgagbR7g+kQX/T+kv3u1e3rCHaCvzkZNfTzzrDda6qq5IAr9JDnDoMWsU4ys39H87Bq1
XPqbrfrQxQqA8scsv47FSRFe6YSfCDhxYXNW41e3BvJpTnuvC8gWD42jJK4qMa9YBWkfVhoEq5PL
Zu1DFVRkgMyIVNRkqOKu7aWQUQ2LL5XGn307C/3ncCz+C4UiUoL+RwL/rbKd5Pid4I6zlAlLI46x
cKSK/xFWxXynqZjP0MFqBlQeoveFRLPnI+ukq8EcAGkzQuqzuv3W4mDopyJMQ/onTCZ1p9YLoBNu
R4i+Fj8jYXDgle0Wra2EwQl6y7WnJRY8xDqfOMEn1vNABseWPXuDfScPDXL0mH3CeMqM73M5b15j
0KlvWBrl7OIZDLZt+Vtaq1Cp6wSp83TWNG+en6ullJHagvfQU3OmyUZLEDsxO4vlIHUsltnQCqiv
ANAUWEfhLRQ2JLTw6WKeySVq4T+HzAekOlfGAPSvgYEh3+GOOKRA0AbDAxeBX2I+lllECR9pvZjQ
oqKETAtvLlqk/50aLjOyFE/z35skwnCdOKq1ACVpidF/wpNSGeM3FrrX8FWK4n7MZiW7F/PRt/1O
vZeh2rghhXrH1EzDcdqpXt7/bECTmxVY5hadbF1iPRKUz7L1qNeoyauHkZRqHkdi1a2k7bZKFpsB
0IveztkhGv7qZ8uS5RNn1xRI7sRiwr5NHWUJlnE9uRLOzpJOAwInQi3OhoyXKRj6AB2hukX1J9U/
pLhTMV8RSIedzNZe+RkzB9hAOjeSlwU83fHphvh5UUj7xqxsUMC3r1fUw4c2bGYwfB4oEVFhD12/
TDyecJNltXHEqC+H/IVUOyLh3oDRoCzXnIDY3rNN9WTyYftpZLHqVdsHJLRD1U540Xoh67OlOf3A
PK2kr5Wj2yH0gDj+2c2WIyLf4EmIaUP0atD5XZGY/UokcO0bhEEZYx0YaPG8sJOqhmmRF1AthYAy
0/tuagrsKqLhQllV0IlfgOdF+h3Sc81VA4JOFG1e73heMaTIT4fod3cxGpAw/jaEqs+1qjtBFbLF
H8dL8XvaaU7zYrenyUaFf0shOCftOPpzwmUqaiLI+cxDquvoSNZ37uqjFhnCPjubdn6TvrCD0wzw
E1+A8F7vPSJjddSb/0TtjqnZlGsm8VVGu4SK3h2fxZ/f1Zz8Tn5AkoFaiZOoZLMGqq1aTFBrQsYn
6/POZhfpFEosa/ARc/IWNC/mCsZYruj9OPaa9ic5Wb8SDvUqRy3eCRc2qQ3AgCAGSzsTQaA7qBXG
lpYtDhW1x7WprgZnshk0L6fDMm1qv97i695+lJXfphkMw3giuzz1xZ5lU4WqK0Nt1wwD/svYq0Qy
KAD8KFi7FV37K6omaj2yj9y165NXSq1R1ghHLUfuoVaajAKjNt4dizE+PDjpuzD2GDJ7NDFGGBuT
ph9QImfyMx699ggtOwPq43RQixl4fM+d0ddevC0x6ciMcjb0hS2CtTPeoy6RflgWcUbPAMQjTPB1
mXtjfj3EYvjYaibzSM6iYhm3CyC+GfUvijwh9NTy1r5V/7OSlZkNCWCF6xLnokPeScADEI5oGEmZ
lOv1zV2p4CagPxSIomBgxN5bolgM4Q0w21uBH0qdICXHPf4vCJg52HntsBcLVzFpXIxbyNGoekPz
RZCBye21PbnljPAVg2TtHOvt9BsyalRx/Gsw6ttp6euQC5PKVkGgu7l4dDV9OkcSZxmIBb6Gmte3
8EMmVNc7mTb9xIPgxYdZl/G6E2/Sle7CcZ61dpW7g5NISO3/SXLKy7aY+uutN25BD/tG/V2JFz7M
/q18ZIsBmXEJIZeTtr//mq+WtJF+FXm1/O01m8dfHVsJXFX+gmt7OOo5BNbwA+dgBL2imflseAjt
kbKMKRvjZwCI/dzRfKJX5KIEJpmeoI4kbADQ5FtXup4C0upPktyRBJKt3iKT6ZWGxXHgHfqoEXnx
chM0RdZLp7DoFzLnUnEpzVEFN/lipOQo9PFg+NEKR2l6TM1kEc4T+hRPC2whh9RZXH9tUOdtApOu
CMPfrijkdn/h7HIOtYSP7+sERmBRmPtGLbK8J6xqj4BwgD/7tmYpbNuEJtXdlCMBEOV/LRPJugHx
7bK3LuPIfPbpzbhYSJWDzr5OYj86Nt0r1x66Y2hCqSJ/CbeyZQksr5FtGSwqgQp9Q1lRz6QmivhM
l4jbROYnCd0lo3+4F566R4bOKSuw/6PXfhDF9cL1IED8Uyv3lGQLk8J9nalEZiFRpqXRB2gYcnXm
vy5evB3qOtjkCE32XWmFeAWSV/qFRIxO6mGHWsRP/fdQd5BR84M+9OJR4pi/5SOmi1bX/ZN1xlNM
J12ibs4wLpZPJT0DV8iQXi0ub1PtO/RTRWIgYMMlwG9t2W390H7r/0sBN4sHeATLRCEePAh2fG0M
ihaJmOmmCOrnUWF3ZfpclA4edzsXGPpjy+0LvRratB6gokKs2z3glu0US2aZhnZCgDobyviYxTVq
aqu9t4uLnA2MDYlS4pLR4zSJ9InhzgkFqp9eEQkyaFnu9LpxDXKXKbQB4Gk+4Jho33Es+eVxiNiw
SBNit3seWnVljYXBg5s7qUgY5IPpcz/spttD85i4uyYX5N6mBfX7qu/tgVYkQteD1astr2EKYIad
mn+fT/MA8b69sxrrt1obDp6N2+ex5d+siafc1TQQDkcZ4QbBZ3WPBnmLz+0yvnb0ZKybIxIdwGPr
nuhBm8Ar80DQhUZrWcWFYD729guh970oXKc4gxSTnzxC4mF0iUV5p4e30vA864BRZcI3fUwbWmv2
toTdWWfnkAOsHFi3KUNLYYegh+jWgDSTOuIgyMlEm11wjRyPcwJ+6Ff77kH/MHgdkp9tqeK0bNq5
0Ss9gVhyQdKaSvSlFwn/hiVXPN8KfChot2dE84hCrCH0nyW9/DqpCQi8kDRokn2dYKkI/cjddFcx
4b++9j+xeMSB44wI13uTyq869mcM3SVyuI8o3rw8MJl0JO6H/zFiORVBexuTFHZ2GPz4CcQ1/rNb
sDlIarJsDmU0Skz6Y7JiHLsfca2qn1vkW5r+2FNiBdzRI8vQhN9srIhXccWRn4FugPZOSd3ByYxZ
DhGtjpbAew8DYtGegCQ9HHgHRUZYjCo1ONGPIVRrpz37OmkynvmSafr1Ub8pwEZKqGBQQGaD5OR4
b89TVWqkbXVRYl+Tcx7OBDWJIXq+2OnYMKUlPV7U2+sDhQm/DQOLstvpPgxDiis2mqRTCYg5FJ5T
3sA6t/eTwQOEmachDckJWHvHwvRfCBtUMS9eRFXD30xUN9OVsP96UGPNj+i9QeNc28KNgcAZhfve
CloOiZ8EHIMpDDmvcYKR8ycHTZKtWIdVkSMqogHmp6RRs89pQaXMsgxqA+M3ScASys2rTRm3Bo47
6/EvaIGL9tGBGbj5flPvtO9F9KEfLNVFy7svrDnD3Nlq3+8z/uz4WxG+Zc6DhRK0MOTh82DtSs4y
fHUu7LvalYXsKEb0NO+0GVQ2oJCxTnPnF1lwZXj1A1Z17IJNRxiCstyZ8MrAiAuPMm6x5ZmxKoZf
+w4OPc/z7IXTmzMGkPpo6T9K/xMkue+HduC3rdwLDrwJBLisEX9Ge4puFLPNK4lJZp/IB67EzVHL
MeWBzd+1PuGfk/LjQPB8cfoNK1q1H5vyzQjD4biYTQ8zYH94c7zo7RC1Atst13f0oLyw2L3GnQSD
f6PnjAZe5U1x4+EY83m8V1sORojoDhdRpykd+YN5HBRPvWQHAIdKgAjh+FLj3e1vHtFk8D9z5YIL
tDpnDFm2bGsUgJJzM1R2NLdm+EAyDgqG1P6Cy+naS0oDBo+lJLJSKBFt3pNv4rI8CmulZpMAtDFq
OpcH2vaLFASlycmLvPAEe1RCYEp3U0wg/8ET4PQKsGRuiOQs5IE4WovUYU94i1m8p5VKv7nJwBm1
Az5PAmPYt4Hg34OKUcAxCu01Ck30sSf7y1KDt7XYJ22Bu3yjfepREsTkr6YRW/kiOTDEwZL5Huh5
TVsh1qYpjCU8LJuYXqPdf2dxgx4HlUv3X/XULPmd5YONUBecY45eVDTWlol5kaWSuA8Kc+UNkYbt
+21YFzdZQIXxAaC35AWflh98Y3rIy5kaonePEwMj0Ljuhop/QfifgEzFCyuZ0Q9cS5cdoPnHWNSw
XqVbk+4uAFwFmn1er2zulFwc7HuQHZpeJd99ZtF6vD3Ms6FDU6UKFd1TxgzyYCPuuKmQ2Pm5tFoS
sY2hzuBBXZE3+tVCn6FdnAGfLVTZW8mXzO8msj2NtOvRI3wOo85nm36v+z7R8wmE+mujaN6sKn0v
CmxWrBkg1MXzEP5nNtB7ZiH3tOUDzHE6vMtajiEbIjr3uTJlI9bTuHtDp/StLxiA1sRv6WFSIRbC
DFuTBoljnU4mQIQUkLsOmsq8b4lJnSGxupbmtbsi1ozir9BztR5kYmYtlhwzMGuB0H5fo9PwPWdC
LDeBkCphSSGEyDfc08cQvnpFnzH5M3t2O1CSixKdEi9a4JrYqmvqpO3c97TfLtfbBv7lfr+9jLqd
VlekZqiFSMgvD+aF6j+ItccCzZYy2lKK8o0zW8NzDOaVBbMhdW7gs4kwdwliJCigMxeEtDIO5UmP
kORvYXUkk/IKWdDWkbvxODbzqBCPqLbqhrBO4S8c7H1KBGQLpv9chCVMBvXSRiKht7j8hqj8MGxe
goiAiA/MM9FqvD3/g9yLNjQuwy9JxOj8dKT23qmIiF3D7kWdwW7g8rtNZGBphRqz0xOhOWfa3YUe
OGNtVv9maXOMRNk8RUkp2quCjNv8glCTa8qtJpZY9gSzp6PND9ASxzCgp+zFp7EfmsDBMni3bchy
N0mK4zJ0Wix9+V+jCJdAZx9QyzjIQqEymajD0Mb9ASKj/onPeAbo4vmgukyiiTex4fQkXZOOEUD+
z0JZtl8LTxLEJ258iGovPOYPYOun9fFvoNEBuxGjI9TUV+WxmDwOeL1G1wkcJR+Fy0UlMmHm3Gpd
AWHPsEVL/L/gnBTdu+jw1FGo9IvQpGlpLWceN3sVAEfVXYQk8J9gpak5Z7NmeE4vJcfIoJGlBdfj
rNh7JL3Nk/Kk0iIRkjY7n3oWorbbknoIQXNWf1qTmIu8khA0xLZBfco4Tr5u5SfhREIsPUpAG0Hb
9Q6Vz85ykUohbwkpVcS4w5LZuCfZkhG6hbBpX3AhHYtABfoVDUEAsJO0RMSapQ/ZFTHAFcdtXFsw
M3sOr1KkNCcTdBcVdvPPgh93cXkj/zGb/tvZ6ikgrMCl6D1xz1SfxtFIFMvPJDmHaRHWY+yS0Kcf
LWB/+EbVp09g8fchojJuOv5+edvjcWgPtFvsIBR+2WF7PAoJAsix4q8bO5cife0zwJ06FnmTV2dq
eslfUkJv0Nvtgl5TB4Dyf+N4sVfP/3UHi06wnTXIfSOf/8+wt68nD6xstcG8p2mQKH9F7KcLP3yy
4QkknwakspWF+8HubDpbMC59LbZbpO3WpEo3cwQb72u/Cofi6p3MpmQtWG+sjh9Vx3LCgN4Vg2He
VTCE0kcpz2mioXYx6yZZ00U9n/aKDwDrpZmpedapk+b3uqBRYrfO/Vl3nk/uZR35EV+0qBFNykPU
N8VBf3aVBXoaq95DpfBNLnrENJoGqiZedpJpmD6VfmMS+Pxcc210uyqf7C2rSkUMK49QrVdN/V0e
Rj0b+l9c2zLB5rw2h+f1AB8a+5MYJPn3asy9pG6VAPUf4b2ZCmeJOwUpaEcwKs5Cyy5R7Er3fNjM
dLzkKOlxRmeRF6B0RwxjJYTJx9mh+rJgLGFdSmg0XuewlR0DlXD8a0OfFF+T5P2Dx0SwPs279Rmr
tvIFXxfv5RXOuhU40Gu/hPsCrNxBnlUJq6ZX8UM8S4h1xDRd3lrJkxowd+UE69Aym1PnyMzvOTWb
EUy//PSz1cAawMKXIq1T+wIaQsUMv9Rkfnwb74Hp52QIgjpyoBJEbZTCr1I56uZUJmeLjwWn/9p1
Z+S0STFm/PQLnPM8suksF4emgr3yB72XweWlKLu4dBUSgk/jLy+L+VrTR2TSt2dDfa8nItYXWNBq
EF3QnVrnLl3dKkHn0dj509U5GcT57kMUCzj7cAhlnWMqbGi4v5AzQl5UqI+Qi6NABUgCIJ7nyxvM
mOJpSB5aCK4KXDAOV8qtPNKZveSQbqGOZIkjfk22ctWxdUoXPgjEWI5z0t4Q5ysI+Zgu/vuMWSaA
LQA5doioasMzNa/iePNZJPVf7roQjN93rMJETAPp1vqRKQq4QUIqu/6Ie6m3t+1RrRasDJ5rETfy
MBHQUijosr+OkaS0TWI0Y93nd3G6U8RIfwlmmiOENokAVOPxr+DLtLdlra6L8C5bMUvpruR8uE/P
oa1vRdva2NsTWgwVLfp5RtvYbTnT3SZM+vV2q3+++gXpi3574i5isBIqPtkk3ptkdVnZGff8Do5p
univhHcyE/7MKhQ/mgMNNQ2n46lr3HLFwcGIypfNgMklsR/G38Uv69VJJ4pPNa02vcjpwb49z4eQ
6KDRoe32AjOaEBKiHfJUgn/1z0AhAWBdK9YMmr4axErvLlOkSUAX1UiddNRVVOysmmn/BdTzU0lQ
1ASdkJCGWoiRs6l8gOK/c1/p4KA7H0BFMaGLURI/AS1jNK+ZxrH4y3fAA/mCSG44a+SS/6Uz2j+/
v9+W4fY3p1ZtlmJ5TaPAEl4HKFK+8Btsu4KyDSU23lhYMvz/c8F7ITGzeRgLsCNc842TmTqMhtGd
EuQ57eSiSRz9M1mVI+rLfxfduzYs7lCF33wgm7PIFXHgH0/ahZHy4e+gwKe9JjRVqWr6djFCWhPh
O3aG/k45KY4+lgg9cw/6X8khfQWOb6LvDPsrG7J0BkH3Q/yOyStf32EZgXdqPMcThV2rAARr/o82
Yl94qBSOEFL8l8M7DYR0CRnGaa9E1eWdcq5g5OfcBsVz6TsgtAUkYVUany5MD+GEPwfVb/nRQxik
nxkPXknNukDDJ3h2R4dOwXpdG3/FavcjcEdu9ys6qR8Aw0NYfBZmY9r211hqehLmbR2gEIgsOR70
3WnAiUx3oU4o9qKorbvUqiJEAdtOsDE4JHbtlut81XuByjy9NUlQZvKipvxu2mgjAHCR0WhWGeMe
WunfSTjReFdF1Kjl4XsaF1CYqcJdZstO5UQJhcCu1yI6eDzpNjldBslTQ79alcDmh12mXEuzpdXL
Lj3crhNkiSS8pdecpS6jb8vPSDDhT6725Hq/dD5T4G9U3tUyVrilxrOh7W7qoQN8FXr3DKIY7CJ6
UbZERr1Iyob62vxGXxo+SVQqzS0a/WGz74xB9Qg77381JGmjTi/8wQofZTvTUdoXa07xJEbukZ9M
GSQ1IcHkHJvi6mf01/9JeheJeGVJTdaOyjFP8pNwY73Ws2fkUb+1RCCtgQejmjvZheoxAtBJS87t
WODK5kDEeLRPgsE7lseBZuDWAMWYFixZMiSRyjcskC2RlVJUiwyTSzA2kKGu5OVIFOFgMe1hlXTt
YBe1cziXTZt619uvTdiOJUAVwwqd3zugN1fgceiVkDSNvzqJOBtwhXfMvU8eGMObDloX0fwiVFS3
Izd46aDJCUdWUVLSvnkvS87SnJM1LiiBOZ3zj78KYVSV2IdAfQbIInSnVQnv2JQ1TT+9A/46aRl6
bl+dnEBahNHNNcAhWu0A9F/4ugW3AAXlq9Yx4V9fOXR0GWLk8RGSYZoiZJi7HvFv/k4Q7eLuru2+
7Pb8ZD6RlolSQZ3sWSVtSOT2Msxwo+0PTcHc4cH2bd54AV+akTG+APKv5Eb7rdXjWOX46k5auUMu
bF+cZc8cbHI3FIdeJLqEF0J4HnWfyz8yLTX/XHjMs2IH8U1Gca/BCAt8l7LT/TrPMAhheCpUUmHC
1GQMhMZqM3EVUu1eB4+JIIwl8MpU0eQNHmCTuyjYeu6EB5U+3KfEZM1qoCqKBHvWYqs55HgGQ79V
4+o08C8Iy2JIs6X6YijLnehg54Iq74HZHe22q85Y/xzPgWeOb0pqlumreHf/CgCpQHG24n436nE8
PfkHJ8rmxjB+EqwHuTtcbQttLQFaWqoB/5x05BpYtO9QUAcgwY3J/u8s5o5iCasOyY/2dVK8tje0
u0uauiQNEg2bADpPK76mGIxGOaYYI+L/ktLI5kZGQXVazcT3t123KiE5HdBtCB4QDn5MTcjEuwrq
HJgIJzHn7t0UUIXzyL0z39a1T+aGPm9vQ/ThSp++pCuPy0MpfwMm6DVd8LQt7Gywl4OKQ2tbUYu0
X4rkxNI6bqCQXyF8cK0EakVkvuhYWt8aTcCfwXIZWFXhwtuaCWeHCm79RpiAimroLVCT5gYfIZ8p
TZyF7yo3rYrmMcfE0RsGmr50h9TfQTOUyzP9LDKiaVVHLiybr6chZ56vFNfMiTt3CxoZX+3Sp4Ot
yvTpeBMiUETIj8/vRDaSIhAZllivwzLpWzk54MEzCwamaqMw/BRjd41w1YN0enqP9bv4Qu676hHC
7YbE+22Sw/QWHUTXBfTRqmuTyygZSqZakXukkdjXfktNwU0DZbge16gmRxLINmx5gh5bgTYrsCvK
5i3KjfFmzp5XGCGxIFOURQMADfQ2ZTR5V0krOcYIkOVsX7/qwn8ZF6nEV/emGmxTWV6SoU9ECmWK
OUSZFrXMHpvFOZB2gER3abCPfsFQ0UTHIuGMaK7x9pxxiaS4bj39nMpHtvW3bU8J9V0ThrZMQyeQ
5FEyK+1cRqVUfpf0uzSl//6KckWlDZHTUKpJlwxYmkFu5Wj3gBErzNJRgI47PxW02g/Duck90rsz
73mfvcXFEl36TJGQXbE6vQZ5Pw629yp196X629b6NBsE8NsXy3l/qTCVX+m6KFMJkJn65tGWsSfG
6MMmIOYRMVxrMfpCLVfGILArFfYOnmvwEVhQBGlRaSlUJ3VmlVJCK8OWfDwASdMNxkWnwbQ0LPkA
Pgh787VG6uQv4+hby6NqYEMHsw+pXGDUbXeQFQiJsJnTvPErpA3d5kOEjjZ4Xn/40i56h2pCaOxH
7CMRPM9Qi9diGmYnWOY5KhyLGaO+G1UuOnBLzSb2R7OHLU9cddAwD8iHoS7u2IPgYY2uzgTKayAS
Ac6b2pER30nmilIkxzjJwi61eKQE7ph7xtrWpFmVWCyo8RDrd+dUV4e15UT0F58hf1+mf6eLwZ/G
5Jm0jjeDsqE3I7QZpoifm1R64tTcSHC8Arpz0IPc1g7ALGorHsbzfuy9ihnVpHFZ1uoAeuH7zuV0
enJfq9fK2G9ia7kQf7paLDDpzFTl5GtEEpCoxR0zNBcz5YiLtOOqBOsa5oAijDrQ99i5ZQc4gCCY
tJHjKoJe49uFeSPaCWFjizpyNhRWNVqC1GvUeLwGwdtVzrS+XGLfK8QtvQl4ARUVza7uZLfLutx3
ND514kD8gFRDPlVMwm/7wBMNoRPTAxxUCcOR6lrDQuS+kGerbu1Lf0B+JPQbrHQMyuF67gImuXZP
9z7GGsWvTMQBMsRu5sAVfU+phtyjFcCZ79SWX+ERJ3RAbT4vSfoaDh6i+MC+AnLJ284Vt9VAftLv
S/susuKHiyLwPEl2CTTD0hvOlRgUWKHtHWXFnNQeicUJMMiwaX4MxAcEYMa6WsWhlIYGlmx9cvlO
Y/30ncuZSHPT/m28AM4jJoGU1SM7Yy/99YmoB4A2EefsltPJNdIbPdFDlMfpfrldYeGb8FOUyEl/
gpA1YHQM5v3tY45ZGKyfVfh5HmgNu3WuCNmHM58rH0DHv62aGqTFw/evxhzCPYZLm+mKw5JQcRPW
dNChy61uBRgz9/KiJMc2F5UIP1LJEX1dDU5SicP4eGrM3/gU+eXZ7X33MD90emzOS7U/XzJr/HcV
CbzG1wEI8D8tJbBo8GKbnqcfwYBLCBevNcQtShn5QHRRmLEu582RBU8TJLQ46v1b4n/vNkaTFk1q
bX7HzRWs5RW2CUODPMeXMEffqKBGnq3imTF9r1l9tyQxG9zSo3CDyRI+gnyaieheTb6X8I+5Hxuu
XIFKf2irX8xPjSN9iYo/msgG9fohnG7ZCCYFOBFZ/RwL9HR6enlkbqbTWjVPodkoHSid9bv9khKL
FZeMtsJDpPGE3lCaeVC/q1o0Hi3uDp2BEaF6Pd2ARwFlU4yDkzPe4uC6kGtRvh4+DDcv9QVXfxiD
8OGtFmCXHerxXFNkJRoGqL+2Y9NpEeWd+vgb4CtqHKYXGUL9nPkwWN9mAdHtrIjItMzzxDilM/k8
AVPmOhXWqftf63M9IXvs0/AR7XL8VuagHm/578Bg9vR/z0NHXiRieRc+BsvBkXexfStU2Rvffxpj
4qJ5nBLJkwUlQbXjlXH9M/HwvK7wbvUV3pQ+nMkC6iVUCY7YubxSt6plMEJzZ2dDjwIOI4aX/xJa
IveaPsUQ5QaVh7HbwUAQebLEyj7eK46U7+b+BHNWYR/gcaxuKA++D0UMaQxiNEaUepRurBhTrfX4
P/BqHvcONWIfCECEHjIoJBNRkxKJEi96IcpiBLPeG2IKJxiCRFJkbhcbAgtQrDjgbtbOFw+I9lJz
HBa1dVVXzISWPSf/QflJxcNxuLKbiWfwlOGQaXn+wC4NUiYojPBaeJ0C9KgaeebcJw7mAylWpkkz
T3EoPqHgmNOO2hSpyaRUIoXjndTtiNgDD27eq7w//fFrZCC5YXmlWEOSlP0iK1nNXJsF/4kgnJdC
bARfrRAe544auJxxtdXVUv6CzM87rj6VPSN2pTqXUIvdtfeJ3nF78SsgNFfgx2bltPdy3rZ7xXSc
6Zqwq3hfDapqrUp0njkiNBFMo6G6nLt0delGR1SEvH6s8iF5nlLJTcpvNDBycUUQ35SRzuIcy2AB
U+WYiJ5yDpMl5Y6MHu+AhQSkoo3deecX/zybsAE/Wk2rtRuxz7EZ3pMZGNuPUSH2vFxFxjcwHNQq
ioQHTNc41P+lBfJxbA3SBpNFlXv04IOUsYLSKg3FigxEY2vVqmxHBSi+0s/OJEaqfyDuddLC9lms
TOkRJ/QCZCPaCqr2q8MKDFosSpkPyqKihZTYBkgcxE6kCI5zcxQAHd9hGGRxsDLaE1/1GPIQyeD3
gsxmbEKvsMtMdyVFmPFYAWd7rA57UN+5SL4Nq3MYcrVRMIR/0Y3Bmr23mIoYZ2v1/K1AAe3r7Bma
TfFS1BPKkqZyPpx1csHKNf0KAxG/Vd/5CXvuZ2uc7Nhebm5+iZQwBc8KHeu0kF0Iy80a9UVU9bLF
HPMVf1AWmgOrBPA8iWem2IaMEaOPhjZWsbTmQX/Gkbd/pDq0acp661tpNQXIBvwdRShNI86Pm0jY
LOhpQMintICLoqTftaIiaVGnNwazbEv3uzXByJPpAK8NxJPf+cAlKsGphHSCFZ+qtCUfjbvPVAxi
hz0H/k7uHgVORbldM6APZ7H9a/Nb4rL+pCV1OJuEaSKchGzc0YtHtjrqRJBs2RwPVr3XTI4vQJDU
5e7Mm70DQQgwcCeGkr7MBZCqL+xNbQ0ACm221uanR7dIHXu8gAjsAHeq1H/vw7FbUxeknqw0FR9N
u49DTnaM1uLFQkOuIfmiFkj/7I1r5gCWdZd+s6AR6yjo9QNohOI6Y2iDgAfz+Kxzh99MuJOnOPA4
D14mz8afVFP3Myuv1uaaCJ9ouFfGUdTQ/wM9LOmOXonmWxb3RUte8VOCykEfRalRvsgB/H/QcYoB
6oHHmIWtX5wenFpIXb+5AhqWSvsAOS3eicX9SFOF3m/VvHvvH+suitTZeJi1HxR8uduIZN4uf8AC
RZCpVWvKT1E7V/edrBY0g/b1aAU7bl5gWirFvvGLnXtbmPKdf+7xds5ffY0muOv3+9hLe1bs9jT+
L6Vpt+lxsxoITbw1H2Gz+c9q/sv8VwiJsGUAJ5ANQhltTNVhuwOMJJXXMnzMGfM1m+8tqQww/inN
wRAuleze+rf2Iww7rGfzPJqcLWOHPwFOxhGWhvA0dPLx0zAWQoRQUgY59GT8J2STGIJ7gtBxnpWB
wRwfSyyRImB0zYQZn8UmVO+YrI/XSEFuXWWHo3h5tBpGdK2GuM2Noq5mmdIqjTURcmGffs9uBUik
aStY3Bodk349Pf37h9/UabDFMihicizkDnUPwIpsFpIN0VNgFmvt72aWKljj6XlSNRm6+oemeswc
SVnf2jGZrVf3dJqkFGb8dORoMyBU5QyGxhDRcle1vR8shA6xGQuUb6WgUW4vzctQp1jewV0WNHgp
C9kXBSgYrrz9OgloVbx17xVBgpRyiRFnfQOd+g2YovMYGg0j1FY/z8WNWrYZWAvNY52qZtrijNPH
K9sT2Ii0WeSYrbs7DZcmaWqDUkiz+AmaATap84c5W99Uw62k/UKAQPwVtCNXSlIC90IT7F5OFLlk
8SRHydrJ7Kci1Uo2l1u4rfQq1qoaIPk9RbW7pMYDdCI03etG6cC3GLQ2SlEuEK3A3bzKok2CnkR3
AqhSaB0ArxMnzebb3gMTk8CUFqQk1Qzy88pGCKgikXn3/IYQXwtKlvAn6uMsLftvvvOscGjBTiUx
4MetbYskpymoCUx1wM38yoRUFzPTEvL+0/s30qxkArve+f0WOQivZBLDV3TMcFAwF/wzpvz27LyS
JeFoBt+tV/5p/0M8prpSoL+cE8YngfR/Z1reKleCvbUJ0e25koZCLrdVPm4ckzOmzj9tQTdwYpsz
2UMAsWkitvPi4eotLMNswv0amYb0p4Z9V8GwR7NkEg6bZltSZJxOGXJedmeKrQ9k6bpU5lXhiC+T
/q876WuPG0C/CqtlSyT0zA/VpB+J24di4lhjyJ/ItvyLF91Iv/vU3rAJm+23SLgtpvg+2C9KrHs6
Q4a8yVE8HKwMjUN+hIkS9N+AdkFXYpgVT7xd25taZ/+nbld7CzHePa7KAYjR3HR6PxaISFJ+Z8vX
RdCZQxSuQF8uHw9BPpFyjZmX3C64AQet0LWWKbRp0QEBnz6SduoTesEWL/lJiTPGoGq8h+ybzBcK
s6rjoh1lfGlDU7cT3W5tvQfgFTUoBu0zQDAm5y2e6xNpYXGleCPIKIW+HlJReeOvx3JtQxdC16tc
igHoA9/D8Q6ZA6d8HRRkO0C1WQoZkgLatX2KkD9C7ShjIKHD6nBpq7E85dAhX8tWLDPI+PpjYdYy
EdlNmle5quFwcVpeoMJt3tKV8RwrCJvIDW4zuW1Asq0IMAnrX0+NVSVtV66zOi3duXkJpMwe3bsu
6Z2QrrdCTYgT/Lx2+DKkh5MCOYwh2gGm5vIweufikGvTqkGGhOLXlBMy4ZreVMuOdrqoiq8gKWJJ
Jj1MlB6Tpqq+TWKi479aN2HfPFvL8+Wl+r+DLdQK61r33y1TDOBafRp2ui35k2rEYxzA5lY6HSgM
/4yvLtvCpdOo4RnIIPjC4jP24VxElcK9ea3OSHiNPSgiT7f4lv2ctlw1IZOk7wX+M7N4hLMRg1bZ
7hTgdOJa0DCJhvjT6fm21lih2YzkV10lIN4qN6b4p7MJWhSr0AiCsHxUGY893AL2/aneftc9jk1I
BqXUpDy/fW9JgotFdnZLNvpB0rh1tHPclN7tVEBrZy9xv7wyF3X4NiYlgaH4jZc9yaxMGKbI11aQ
zPzWOLfQsn8ISnB84bTuAhW8kWf89w4igkXkoovgcaSjEiQBb22mCIS9ZsnR2XD7qlTcyQQ7Svxs
gqCoI2y0hxfsKdIhNaOCKqWx3+ng6EHYJuPLpBEbaut0KP2DlAiL9PcQNLm1arI4JqvKb+9xdyv6
/HV7mpB0xO84xWqr+zwJ5dH1P+wVnZQRhvqkVHVsMgUknOjTDYUIrQ/rLEOvEbI5gDso6mW2Jdzs
heDd9AJbh98V58lPrEDK0DGqoFW9/3FacwrBFj2eKKNQIRiFIXeisXuaoNRxa/YKA8RYfsvg/vm2
U5nmfJlX84FxmGeO/zcbEgM1XgYfMbkNT9tXMTf4PtHGLTXHoOjr90hFMnpiUxsy2cgPd7T0Gu/j
/rosvo4Fv7vb/Zgzaowgh3sC48Mu+JrsHvVXI9yb1HVd4DB08ew5Yxo3PubvwbtFNs4jap9j/rf8
ou0EEZZrd3enYLY7wUTWMLGMTIeLIhfky7qPZZJ1aV2qfZO99xz9RFtzxaP8ODnBC0PG4G8dRW9S
SdGxJETV10rWJy+yTT6bU/afbKq33LgmSmlEtwr8eapIA4qrzp1TN/WVbNVvZ/dRjZsrxK9H5f8y
GSZWW75nafiH+oZHkQrjNlNpfxxrOCugjPQ7DqsAQ15jS2EHZCA8D/Hcpd9Tw/NnXla6NnNPo2/y
yy0CkPMswQjlV9CSUxe+dtsjWP79mEsWhqNYAgYqojWN/fwGh4UZvTckhnVgYO+NeM04tYWx5Dh1
KpIsQ/utPO/GqlTB7mB5ppIUkL1auQx0AsbpwsQrwLEzpcpyp3+JDAgdzHQoCKrXOMtlJmR97LCb
HedfJtM3O8PFveXpI9FAzk2bI1yuK0r9NqEtHnyFs/IrfqYRtM/A/R/R4y3/kKhJKPJglxqVIpXM
BN5kIFD3ZI1AW5/KtrhMpnFDTbIZhy8RJgwREHWTbc2jXM+PPz5UTJ+0JFFSAPDyyhIVzRvjUMTD
o4c2mCaYCi9HgK9O1Hi5whsSz774iTAw9LZso19vzGx62GFEvTKMFiCuc7DGWMH7sGxN7HznorPK
huqLZsqHHCOOH5SIWEa5Ia1nNYuRtJNi8g34ao9YgUxoLw9pIJZbtSuVqS+Kjnh4SYJ6ULMrtBz1
AgVlqWGOxgBFXvVSCv1uJ/6BkvOzJuA6/KFW03aqMGg9LlWgYmZTqHj7iFcCBXviKSCcLTBudauN
F5Dny0PEzdicFcL/l82QozQu7U6j/USsiptkrYa6q0ZzSUoPaID5JSUerd2C9cOuD8y+ICBLNOQN
uiSHRxLaFoYbSw6MaOgS014cy8GrN4veQ39ljwz+6+el8jXaYyESGssPJ0jY43P0ZDN4mrc/Ww+Q
j3j+rzb0zgR/ajMV0l8gZQLC+2Gf++ExrKPkHDSIEk/RSGSGQ1iCB6oQrNuwTEE7Brt3cMoN0lin
Xq+DLPhUBPKmWkGWbTHTu3j3Idx22qY2/uiCL93wpF+z844LfHI+UJoFwKAqtARAZ20eLZDpIirm
Ds6vM3hR6HurqTGKkTTOmTUQaaXJYVxAef2FxffSgHI73hKJPit44JNYdf5DDSwyY0zEgHoOilYy
uNF7VyLjorOIfve3XU+6iiTR8TK8H7LAovFZSJyLjo2IaeNkK8SvnynnOv5jZ8QQ0rEfjpzKW9xl
S3i7pSYzDQjpAOHQTYmK79SHe9RKVRZdl80oHz9r17utJpwTLlgti7jiYDJDGwpemoCzXozcH53s
eTNiS8mm6Hc98u+3fpK5C39kjgdEFmzyGKhohFD0XWzzB/vGxHXK5+ww9OPR0RXY8SyXvnMhgokS
VheFxO070U+P7L6dykgYb5vVf41FDFbtj1XmDCliEZWUUVkBNavNiBvEDa4Zdnid7MNxzEYil1ge
2FUzjIk5WXJM/vLqQSw02FonvG9WQs3RRAAreoTmQYjHUPSCJAnFsFaIAMpUqWHVTMqkoKw2pvU1
5W8PYk8p9FB8Iw7hRBMwFrE3qwoZZQRvGYV5GM7QbkBDnPGSEZkLs+euUSYABxiKH4nG4eaBS3rR
BJCmSpWaTMrBE9Bfl8ghgJ+bhKJ/rmvGu72VQf0d4IltjXw2N5xrR23tVcYz5ojHzeZzPMhnYkr1
aLDxIk51ob2rK59vl1WLjiG9QafuymlrlmHXtwGijNotGDDP1AOXZ5sUhpKevoWxk5l62VylB7Gf
PBuZpxJcuj6hteKR4ofBFTUnjrT+fi7suZ9YJBBYq6/2llALln5vk6ydL0pJKhp6rZWFgsvN2JBc
c9PE3c9Um05Lxqs9Rq1DDsQfBwq2gZk8sYSnB6+2BWOyPbbF5VvQbxjz4N6THQJoCbMWWU+op4bJ
xkCrcIu7K9ZpvW6GLBSt3wHckr4SNNUAtaBhCJYRN7BARtB/lUtaSVMmaADste9srb7bVwyoFW3+
WyjsFSzc10j8iYTJo/Pchu+br10JvL8+hn5eYvM0L47L4MlVpxsqcGJ16VSweVRL4A6ClXkovYc3
DMW8kPB2FTDkCY9iwT/E1BNpz03Eq6u07dAZ7vpUQZz/2XWEzpnwYncVgwgQPwAqMa4c03VmINCz
+MvkRLbpO4RS2LuFJ6Uqqa0mUy6XBK87QFgnO78kRlCD1/liXrMHcTlaZIN9ttjZ0ylozBj1r0Wy
t3NFNBfw621eLuAtdHKSwSXK6lyaZey5UvDQCcn/YEyTJj80mV4G2WOhc0Lj1EmSZj24zWi9KHKv
XGgpm0DjcqngW5e+Kzaa7+61KeEwTsHd1JNHRbDtmwteUBhaXnExeQq8tklJKU/0ADjMLdC+wWOR
5LpSvTE2HlfZR9A55U/4oEduwu9jtXAbUQFkfY1+dkcoJP1pQ/P/qoMcKQgly3R68mb+t5+drmFu
J/WHci5ijNARnPN9KRZDgS1HA8lq1zB+MIk1yhjdftJJz2KTNQGZpaHANgKBId6IHFHCU96SAJP2
8F+gpTvKgB9U8MnDIw8Ticf6EYblg7cPfGQqektsXMPCxloM42IvKD6eXq5NqKOd3CrPpTEwb7PM
eLaWN4Ykv4IbOS+BXbHxr/YaTeSz3hEHFCBYSS7wmfswP+Tx45NS8N2AhO3qyhO4qZNS+Uv5qjpk
2dHAKsAAXFhhd0SibtwHMv4MUwbTXeoSxl+af6IcIniy7OU4R7cTKOvWHeunFANdclArjSyWPP5v
rzBcOaIz8dhw24vlD1noxkPdZ1zuhK7p2y5w1MF7HfOLzkBa5Iby9w93w35+HhE9dAWCMnIcg4uB
6jxBAQ1u5Tz0QemC2VUg4DYnDCOPIPD5QoH8arW5X6X+5IiC7iLYADT6e+b8sfANI9I7u9Ddqj2U
gDdFmPrqG4q9bRFcSb0RxoOb8ZGKy37pmgSbICZ9TmcMxjwRVgnxVOCGGxyWL5qIkYV3BWuo/O3P
Zs2MzrMFEAFR8EwmmjHFP24vL3zs9Y0fXeNwtB4sdXspapsK1seIhxwR1iVuWPQ02LBrLuvuKRe9
7TQpDkITwUYz3dWVt7uY41ueKUZKRKq0keur/KjAgbpu8DXR0V1Bz74oiQjw9NuiCzg74APnwvpg
JQ+LyVkEd6uLBpUwQgdC3zr6d3lVqhcjNm//XjUoR31iheXfZduqfPfpLdaiS7xQz0V+1RUIUMxt
nJvQXxLcq201Bd8am+qzliSD1U9QSpPUh1yqcjHj9e+FDNGYWUXMViC0+dk1YPq5T8/9T2CMNRik
By1OE1MdbYbD5GcB283q00P7ZqIu2XpbkdzNiu/OnRqQa1E+OnYq58CCuHNnub7+WIdCwAcHl/jw
StklqJR1rcjn/LSZCTEyXuHyfUdP4Vgr87YeBEiO8ixCPWA7l+uWv/SnpnQo6N7qypgkXxf+/Xsx
lDXJZEVNBjzlFOnP85T1xKNn/V8zF3hszRQXm8ilxfc5Vp4QVcL0YSZPNrVVQIxeWB4taVyv0OHj
wN6vRAyRvz9Piigum+Ds1gv6FBfkQpYByqee+pZ+gHLEGOmyolZs3LBtBpa/Z3vavc/lt2dJk9IR
hxmC9kV6QV+Kevk6DzCK1axrQCQP3sghavdOGYPqAxsNqeHnKxlqbDv4AeXmkkQk/6FDCvEpf5B5
N/LsX9QhpZVvoaCnj72hD9WA4JwBrKEICfWxw1PGc3HuJ3i5sByVtgxHpsgXoohw5yYQGaUUZFDV
GPTA5hTQ2SE81OzjpgNV1A1koMigchDDIedKlZCwLIMHF5UP9isKe4kMVXqXRRrkcgjsvoIxcNBI
vr+GVOSkcHEI0h+G3SuHbMz26QL1ARPUZq7dN5dOlHMiVkvL5uKX4sD+WVhJpyHATDnN5ExYdOBg
lFlc75KD22aS5e/aB2tQBJRNVEWVLPOOJxqiInph81BEotOHJg5NsQdmmrJdc4+xSGh0M+GXD/7/
SvtdcW8mg2YRIP1GPZy1sSoBkrJN4A/7hTGt4Oqn9kcC00/XYZuK9KPob1Zc84aWSrUyJw1UtlG+
ZYGM3bizDw/GPXv+Os2EIZ0+mvprflM87a26/GT4DLxLCYupg4LZp/73Ibt01jwOT2cr0emGPlBm
LzG4OFmdO7IBYcwMJ+fFooHdYibcWCmtkkVlFAYhb7481uzMlnS3kHPwJI87IJJT0miZQBWlYrvB
H3vVmzfcLuRr4U/iPsgb/fPMy+F3kCCWDczjgmizLxfPPZvh0WkeOWlvZH9SWKwK/DJ2STqT1TTa
ZdOalmA3lI+DUcIxn1IyZ4HFaTIOlHqGOHu4fHKZlOeQRU3d/xI/U7mx7QdhYNwooWfXPs00mBhg
o0tQR2mPYYEenHfJtusTUKXEK5h6BqzTfGRKtsCEYiZFjGZCmPzWyoam71bX4u4XRR409C3Bn1m9
Mt5kGdLadzxzanvmV6AyU+LJt3m7J04ZXT20KMFzsBxMIZQEAhyf9E4w/8oDuTB61qfZYg1TV5fL
mppJjZMovFtXcO4czzL4jC4+93012n5TF/N50764DtbTkr5L//VaBdp7IRUsCs4jvB3OLmWs6vQs
2YVlZBQZWOAZGyP6Y4rIDu8PcH6P0CNR7BVyfJ7BcwNpMTl9nlU6Vwsnisz/d1ZIkN6RnDx1DSqp
5HzdU9EY9o/blQ38blzN9l9LeeUDGdTop2IiMil7haHu
`pragma protect end_protected
