`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
L0mCJ2SrALU+B1sL7EZNSb6Q//NUmXqQTnC9/p4Ba3xqUohP+sQm3uKmvuOqOn2MyhsNtUKNIcb4
v4wh4afRcg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
IsS7zFob9ooEO3sdOw1AQZnKu7ttt6G70bS+r5aTIF+o/gEAw7m+u95V+M4cqUQwj7O+a/B/Xp5K
0+qKSxE9rmT3UwRzPvt8jAdu8AR5wqv8G7QqSm3bExe0gp6yTJOaDj62tyOREvKJoBNnmbFGKvOY
diLfCXIyyp16LogGMoI=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
k+VHcNoI1yKBbiNfxFJ3ERUkIEI7qMJivGSVwlw/lK8NzD6gjhNAXqjmOvn6UTVOoz/wA9NjFkDK
NDWMRRHmtwh7y49atogCtYNP+G6D3nKK/i1BxIgzsXZpz+2CkGe5VEQgkWawuckKTOFrnRhffCzJ
AKDb/VTSAeaILCtC9wej7qsf2Hgb3rHzOhpJ0KTAczTtuVhQCzO2rh4rWvmJZsCIxczmoomp5SJM
wHrt7ddXgJMOPEToaE81eLnQuOLBaF53L4ZiJTCZoQwaRscjVKq/M0kSyOq0gzhQEIRAxxL1ErfP
hGXBSFoVKmlsZn8L5SIWWo/ZSiySOoNXNWe2Mw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kMBkgodNiEQarNwSHS5T3m1CRazUra0Gad03R/MsMVpnBTPaKwoFCTaoXK/5lPJUqo5ZmU4jNPIV
yiNEFpp4e7k6FWDYIe2LnkWPfnrb31RaBoR107t4b4X7P5h0p+cVPcGEBsytNCOGG2YXYXhuXGqb
Yin2H9Uz2OlF8GvpnZNmNLJDPcQzoCw9SZtq58y60zAGOzlVRAczcrzQHrBYpZTwNo4SRe4LHttu
ctyadd52G+xRp/eGxOxDJD3WqAee5y/jsjKUp+U0GECLCZvjQeokvq8C6PjAoPwnBLtMkBd/gyfT
GjWYBYXvxLTFozBmfS3ECdJxeXMn7quR7iECDA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
rEqVI+n/KMvr9Oq1xazuhp7p33ElzeCKyWpnITj21NHe/e/Odo3eqwWQBpWS5VYOK5bJcpkgyQkK
xm1LbRGzVWhow+OLK3xwra1i2Oy71ulmjxIQd2b1befRpE7yOF6LAX53By0tdvsyQtV7ZTl1klP4
vRUh7FCR2N2CTKCEynSh0oZ2jFx/9Q546G+IjC9OJGT9iQ0iFt4tAjLqEd9Svp5TyugkiGGF8v2T
ymTFY+ncTySewyXBFCEw7GPh39m/CA6SZgF4SJGMzgYa+A+O1UJ1e5f2Cb3soZANvs0CztcOOP2a
hLNDfL229SQGrigGWsiVuQxsd0/MdwraiYRlRQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
enbB4lEuxurzSV324UPvTsiO2jAosYntVazxHN8a35h0eLRaGXMlOtluwaSGcdlpvQ4O6bxogVgJ
JoqkRtOUJY0Nn7Y2eMtwypOGxBS/kJM9821Vni3TbMZAR6JmQScH+dW1lkUDYDWTMK4hNliJVGFq
0pkVgn6f7q+o91zVBvg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lYR2TpcVRp59o7iIehjPJBJvgBkpyv4WkukTZmZu7Ri9cNasODRNo0OfKnDPJBytSiKE4Px9gELk
wy6XtRYOnsUbURO4rfnLlP2UGDX6DzxRPMTGxI79betJniUtDvZ0NkGo6KobMgLZQ4mBpAcP+D6y
GHeJKtg6vt+V5fV7LejFTbT5RqOMoGHzt28aHd2zxSZmBQTj1XTETmP06byQLUT/ytGT3qUoqhmh
2jE9g8dhDkJF2095uEFBwjfSDqrl1ttnly6xJVBT5tl4MShkUnMIDcJ/VJvjVWw8noU3d1st0LJj
zdEz9bb9bOI6dMru9gZ+IffHr9M3TKR7k3etjw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3136)
`pragma protect data_block
AqU0l6/9QEVFIhNL0JK0DeHM2kLIaLTdi9w+vEEsN7xYLJ/qmeW8UaGVKttRcQ7ifw03f08IwapP
pYKyFdDE3TjCwcjcuafqmmRwsUjAqaFpGEGjkCIhVxgREtmb09KbOxMuqAFfLgBXJL0EEyd9cob6
l+8W5RurbMaevyKE5krNzGK4MJYZzToScHFLAputAGZMK7BH+v2VgTzsIvjFvfbMiYoWbazNIyYj
k4BQ3OGV5PmZsNbnH1u/B60YOXS2y41dFldwQaOni0ctca827rabRnSI0cNHVn5eC12JD8+MWcdI
PrKa+PUr5bIvwQRrexvmz0wXxZdjX/K+UR4mkvCf3xP4ADSZabqU0YnybFY0fYOj9hK6K+wkCkCi
KyUumUw6K9I+WLlwIapIJPcgHvQ0BgdnxydnfS7soyEUjWoLxBXuGbgDJBWtJ4lFDGgOL6RMqIU0
MS/PTiWGpuU4eqmydyWGEAZd0PRYYXDk6qTLXA9Lqgtyu3i504qP4KjYMEqFnJBfZB3V7JxncuKI
TWdctlN9beyXxtli2zVhdJMM6BmOb02CJ8EmII6peTEi6N+TOvIDzaSN8KyZI7BH1Bcrqb2bvySW
M9M65ZNTASpQ2xzms+yrR2rpTwcxQAuysCRCUpbX0n+U0gQm5x3R/cel5i+cgCHOArk2efsa7q9Z
s4r5kVkbAOZYNA4GSEZgZHuC3LxDYC+TE7ke2Ed0AWbWtD645eeFcc2GwQ0cjz5lkNaMQ284PuxF
WgY5o5VScp56nh2qKFL7Hg9HBmhskeNwBWId0Bnv0pLSmV64i74tNXugXDt50eXCalduw/1s6TG8
A2qnmy3tOaoZTi7kIjGwMLpE0My2BnkUJ3CoJOINtRft32REnZ22NNTyH5uwNIudcBTs6/uX03bP
qC5KX4x1s+LpUfGPdhdoYHmT5ZVg4UgmB475ePfYieTq8vaBEQGntmCpqDKK8ju3E6PBFAJTssBl
SbMXzJp4o7DU3vbw8dZBENA11B+uuJagvCo4PnUSG121hc077/RR+uP1oSax+2aqhrn9rUchCrho
EkFd8oGer5o8Ado6YZxePCu5RYao7qeGQvOsTf3/My04GwAVSA3gYNDpEl+JG7qNA4sLYv1oO9eT
X96EWKoVeF3PT8tEFOBqDdnzROR2MR5Hq8pvaX1JiNt34DBhtk1aVczclfFafamqNQ/wEyCVYyyS
NoSYWrQrtQyiy7DUc3H/R6ANFxCo1DO5Ffs92fbCT7yjxJX1p/WBBNnCdKLLzyJb8iEQHKieb+o0
6oFD5xy4zRfw29G3dSSskRj6fUd7a2scWT0jHcUB4JSmoQddGlDkLPgEwkeuXPMdJAJ1D1pxcq+Y
GgL7+sLQTbhpAqqnwzicWwhXhd/RWu7xetY9ESwVkvGA50sOgQqk6xI7iRv6umj/4r2K6SOlcyTs
MgpVXU5DNyzgIKZKXM2M72EIigegTJXZnEyu4AIyC3iptOAFWOkT69RiRpOUjiQXEVqtCXEas/7y
xOW6xA77wNK05e0t+v6KIpqL/xFbOMMLrnIUkM3OzsHZVwnYFKSaHGeKfNJXWPU8t3h2kBeJGZOh
LozMAfr9MVa3moQ2H+PD3bRiCmN1pz45k5ELQtNBxp05puOnPVw+TNJB3l6QI67AB879lzhbz7R5
NDsc4+Mg9Gk+MZ2VIYMqpg6OUd7ZPFTvOTIwj3rwmcsK6H3drYX5/QY7XsZPWjq8fLq0dCTg0nBZ
VP+GBUeTrxOD4yWrwJCdNcvzXlwZueO0ho0SUnXX3fWpUW390kYZyFZTGdEHEVjorCS0XDnJSCu1
A11sRV/C2xVTZ/vXk7ahquv5U7TYwObWkuoW/FIDKubHGGGhU4PcX/XT1KxeI0neYPZS22a/w1K5
dwZT+z89uIeRNCshY+VW2ao3KRgJ/uAcNGT6xlzepxiFJik0og93EtuADnxvOPXIhuAM7/lxCzPE
EY6gdj1lbj/vGif/1F29qMXrGzsMUSHBzwhhAOLTw5k22CdJymE+wXjgdBTWniXgYanOXEq+/mns
N/MdyZ+40n/drhF4HREUQ4oulM3urcll09Tich2h5PcB016oCAyk0E68QO9Yuw3QV2nB2QUZ3lGh
lT9RYU+2UBV0GUfUaWEjPp2AmVagCvarj8d8DWQl3mlDcpanEz9yCx1a78Yu9qLmaiIlne8qajF5
HD1UEZWrazrUYQmTBQZorxGO37w5T682XgBuAb0uHUip94w4r0/XvvQmPF9BB2OCGcyYLiv4RqAl
pk9nxC80iVunyBz0842PvBfsrCTCYbagBvamG6mwFH7VgXecLyjkTWFmDc7j9PqXJSAegm72F0Xd
KtFpg96N/Xe8uWwgBgNNeBv+wXVcs6mflTxOfn00cIlHWWJ2+QKb5uVPhWHL7lpSiem3LTLVyUpQ
rc4UIZPNlhxukDn2zVV52XdWhj8SBZ1PCBpjWAdbN9hFaDu/2vGuXYFnW/GLIGHOiwSDc+moif9w
f/Dwq3VfFgdJ/cM2iDg1JfkxhgCesZm/Jr5Uu2l/TKrupZgfMGyrmLSbVFEgg790rhgj/nTrJmST
v6Ixnnb7N0q8/JITEjSuU8AnLwimTQlYWwEg0at1AtWfhduKYdt7pw8NFhEt5Tb8Vaw1w/Nd+5aM
rQ3pgQEE2NHjShtQTu7fP98SNMphHwa02l28Yz7Rv5q+EqEt88NtczK6C/GotAuzsKTfgZnQbeuJ
+XU2k2wRIq2kKWFtZFpt3lov6jI5DNg71cl+r2cIAIX26Ql3ReXCr5HVOX648+su5ySQzQWZ+ywL
SO67Gjc3Pz9mG3+up45Yj53hdhe8yAu3K0h0GkOIB6moJULt9c8sd5NTrYBvsa/uDEKsJVV+soq2
1hDWnCJ7NzONe6bXbl/FN891E78BijTiggEU1qRVusTK5ndiysZ5UpvaGg220pjCZyUMazlwPbYS
okoRvOrVzTWWmOVoC4Myu/cCOA74zyqqrJ8KMTMfhpTExqFa7aaPxt+JkoHV9k7dzW13BCQf5R+V
AvF1bdDEgO4LyQlsGhhrs4vNBIHEl7F1GI6J94K22jT1u1zouVzvn0awMCgXuZOBF0DSlWNH3XqO
PKhnuRJSgMnOoSf3zsqroF1YY30cQqzWDSEAA6F+0/N7E03f6KrDSR1+zyJP45/dM9XASg1HRMLR
gsgDlXzNIPV4avBDqmy+KMhP07SyUe/FunyVPKIBmyXX8W7wMHqe7pndSgRySVyotmI1REZl5eqB
YRQtXDmxmaowTs0Bc10MIh6Zs2/eJb+rDVRuzTXIfS8lzcg6xzLt0fxN4QwAcwV/J7uxEWSSvaQw
3es+x01bcxV0cTk4da9l7myddCoAVLo25CqULTq2P3qydjd+lKr4jYpm8pj5JSdkc4DQyIVn8fta
Qyt1KSTgI57DKDu4HCSqUeK8nrmW0w5aYz8Pon9vAgt0rcLVLjGdRsq9oekmhOOh9iG1SYL/tjD3
NAjBMaB+xk9yRKAiX6rg82Xxy+yO3SPUHAJJor9yFJgV+SzNWB4G40fYuRFwFS8I2QXeuf0Sy5TR
eZUKBNnEO2/x/xz1iQNjRJHPnXX69f9RitwCnyaadhJVvwOA8AhBAtpB/55/o+seKDJYL3fj3Iiy
SJgyXZquqFig32IpbaJRhcrukZ9XfXyC18nkiPGrNeh3uCwCFdgsOiFVitOy4vJcvmX1iftQOKIz
oLDRargHwJrzggyR1GGzBhU0/oWxaQHA+B9lCnAyco1pIGZKXtDq2u7hO5h30rwArj9RAaQNFQZL
3NwCAZ2rf10BgAJ5FJ7uvsmCHHYrpiyzkmzo8OlfJz6+bfyTcK+d8x9fhXhzsgHSXWXekl4Szls0
FvEQH9h86XwaeZkcSCv04W3Hs+RBX+rLZqUg73I7hWXuKpX2QdS9GUxfp3gfsIeIgy1VxM6R0QwD
IDGATxYObvguhZELcpOFsyght5vHrmV85tEeswk9kQb8ZQ+MT+vrT9BJHxWRttdjVb+qOnoBzvea
ioRjCHtvSjSmZ4XAdPhKT7DPuO4sB5OlqGt4BP1SRM5qsiHo4At+RkztXaMbH/BkkrKye2KySOPQ
QytpwUUL2jnJMuQlJWU0Sw6JtDSryxpgMeYUTVQq3UTLDSmyh8gjOZWiNjd22QRIqp+uWT4C2TQH
BA==
`pragma protect end_protected
